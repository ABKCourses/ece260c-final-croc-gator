VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO core_wrap
  FOREIGN core_wrap 0 0 ;
  CLASS BLOCK ;
  SIZE 674.88 BY 700 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
  END VSS
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  2.78 0 2.98 0.72 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  660.38 699.28 660.58 700 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  350.78 699.28 350.98 700 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  353.18 699.28 353.38 700 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  237.98 699.28 238.18 700 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  355.58 699.28 355.78 700 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  357.98 699.28 358.18 700 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  360.38 699.28 360.58 700 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  345.98 699.28 346.18 700 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  235.58 699.28 235.78 700 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  365.18 699.28 365.38 700 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  5.18 0 5.38 0.72 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  367.58 699.28 367.78 700 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  343.58 699.28 343.78 700 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  369.98 699.28 370.18 700 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  233.18 699.28 233.38 700 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  374.78 699.28 374.98 700 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  341.18 699.28 341.38 700 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  377.18 699.28 377.38 700 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  379.58 699.28 379.78 700 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  230.78 699.28 230.98 700 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  338.78 699.28 338.98 700 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  7.58 0 7.78 0.72 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  384.38 699.28 384.58 700 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  386.78 699.28 386.98 700 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  9.98 0 10.18 0.72 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  12.38 0 12.58 0.72 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  14.78 0 14.98 0.72 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  17.18 0 17.38 0.72 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  19.58 0 19.78 0.72 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  389.18 699.28 389.38 700 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  228.38 699.28 228.58 700 ;
    END
  END boot_addr_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  391.58 699.28 391.78 700 ;
    END
  END clk_i
  PIN core_busy_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  393.98 699.28 394.18 700 ;
    END
  END core_busy_o
  PIN data_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  21.98 0 22.18 0.72 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  24.38 0 24.58 0.72 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  26.78 0 26.98 0.72 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  29.18 0 29.38 0.72 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  31.58 0 31.78 0.72 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  33.98 0 34.18 0.72 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  36.38 0 36.58 0.72 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  38.78 0 38.98 0.72 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  41.18 0 41.38 0.72 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  43.58 0 43.78 0.72 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  45.98 0 46.18 0.72 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  48.38 0 48.58 0.72 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  50.78 0 50.98 0.72 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  53.18 0 53.38 0.72 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  55.58 0 55.78 0.72 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  57.98 0 58.18 0.72 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  60.38 0 60.58 0.72 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  62.78 0 62.98 0.72 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  65.18 0 65.38 0.72 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  67.58 0 67.78 0.72 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  69.98 0 70.18 0.72 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  72.38 0 72.58 0.72 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  74.78 0 74.98 0.72 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  77.18 0 77.38 0.72 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  79.58 0 79.78 0.72 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  81.98 0 82.18 0.72 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  84.38 0 84.58 0.72 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  86.78 0 86.98 0.72 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  89.18 0 89.38 0.72 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  91.58 0 91.78 0.72 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  93.98 0 94.18 0.72 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  96.38 0 96.58 0.72 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  396.38 699.28 396.58 700 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  333.98 699.28 334.18 700 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  225.98 699.28 226.18 700 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  401.18 699.28 401.38 700 ;
    END
  END data_be_o[3]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  403.58 699.28 403.78 700 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  331.58 699.28 331.78 700 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  405.98 699.28 406.18 700 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  223.58 699.28 223.78 700 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  410.78 699.28 410.98 700 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  329.18 699.28 329.38 700 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  413.18 699.28 413.38 700 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  415.58 699.28 415.78 700 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  221.18 699.28 221.38 700 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  326.78 699.28 326.98 700 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  420.38 699.28 420.58 700 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  422.78 699.28 422.98 700 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  425.18 699.28 425.38 700 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  218.78 699.28 218.98 700 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  427.58 699.28 427.78 700 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  429.98 699.28 430.18 700 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  432.38 699.28 432.58 700 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  321.98 699.28 322.18 700 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  434.78 699.28 434.98 700 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  437.18 699.28 437.38 700 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  439.58 699.28 439.78 700 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  319.58 699.28 319.78 700 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  441.98 699.28 442.18 700 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  444.38 699.28 444.58 700 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  446.78 699.28 446.98 700 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  317.18 699.28 317.38 700 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  449.18 699.28 449.38 700 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  451.58 699.28 451.78 700 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  453.98 699.28 454.18 700 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  314.78 699.28 314.98 700 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  456.38 699.28 456.58 700 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  458.78 699.28 458.98 700 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  461.18 699.28 461.38 700 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  312.38 699.28 312.58 700 ;
    END
  END data_rdata_i[9]
  PIN data_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  463.58 699.28 463.78 700 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  465.98 699.28 466.18 700 ;
    END
  END data_rvalid_i
  PIN data_wdata_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  468.38 699.28 468.58 700 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  309.98 699.28 310.18 700 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  470.78 699.28 470.98 700 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  473.18 699.28 473.38 700 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  475.58 699.28 475.78 700 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  307.58 699.28 307.78 700 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  477.98 699.28 478.18 700 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  480.38 699.28 480.58 700 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  482.78 699.28 482.98 700 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  305.18 699.28 305.38 700 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  485.18 699.28 485.38 700 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  487.58 699.28 487.78 700 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  489.98 699.28 490.18 700 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  302.78 699.28 302.98 700 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  492.38 699.28 492.58 700 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  494.78 699.28 494.98 700 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  497.18 699.28 497.38 700 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  300.38 699.28 300.58 700 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  499.58 699.28 499.78 700 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  501.98 699.28 502.18 700 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  504.38 699.28 504.58 700 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  297.98 699.28 298.18 700 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  506.78 699.28 506.98 700 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  509.18 699.28 509.38 700 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  511.58 699.28 511.78 700 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  295.58 699.28 295.78 700 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  513.98 699.28 514.18 700 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  516.38 699.28 516.58 700 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  518.78 699.28 518.98 700 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  293.18 699.28 293.38 700 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  521.18 699.28 521.38 700 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  523.58 699.28 523.78 700 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  98.78 0 98.98 0.72 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  525.98 699.28 526.18 700 ;
    END
  END debug_req_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  290.78 699.28 290.98 700 ;
    END
  END fetch_enable_i
  PIN instr_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  101.18 0 101.38 0.72 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  103.58 0 103.78 0.72 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  528.38 699.28 528.58 700 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  530.78 699.28 530.98 700 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  533.18 699.28 533.38 700 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  288.38 699.28 288.58 700 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  535.58 699.28 535.78 700 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  537.98 699.28 538.18 700 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  417.98 699.28 418.18 700 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  285.98 699.28 286.18 700 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  540.38 699.28 540.58 700 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  408.38 699.28 408.58 700 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  542.78 699.28 542.98 700 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  283.58 699.28 283.78 700 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  398.78 699.28 398.98 700 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  545.18 699.28 545.38 700 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  547.58 699.28 547.78 700 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  281.18 699.28 281.38 700 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  381.98 699.28 382.18 700 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  549.98 699.28 550.18 700 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  372.38 699.28 372.58 700 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  278.78 699.28 278.98 700 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  552.38 699.28 552.58 700 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  362.78 699.28 362.98 700 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  554.78 699.28 554.98 700 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  276.38 699.28 276.58 700 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  557.18 699.28 557.38 700 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  559.58 699.28 559.78 700 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  348.38 699.28 348.58 700 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  273.98 699.28 274.18 700 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  561.98 699.28 562.18 700 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  564.38 699.28 564.58 700 ;
    END
  END instr_addr_o[9]
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  566.78 699.28 566.98 700 ;
    END
  END instr_err_i
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  271.58 699.28 271.78 700 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  569.18 699.28 569.38 700 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  571.58 699.28 571.78 700 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  573.98 699.28 574.18 700 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  269.18 699.28 269.38 700 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  576.38 699.28 576.58 700 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  578.78 699.28 578.98 700 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  581.18 699.28 581.38 700 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  266.78 699.28 266.98 700 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  583.58 699.28 583.78 700 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  585.98 699.28 586.18 700 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  588.38 699.28 588.58 700 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  264.38 699.28 264.58 700 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  590.78 699.28 590.98 700 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  593.18 699.28 593.38 700 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  595.58 699.28 595.78 700 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  261.98 699.28 262.18 700 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  597.98 699.28 598.18 700 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  336.38 699.28 336.58 700 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  600.38 699.28 600.58 700 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  259.58 699.28 259.78 700 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  602.78 699.28 602.98 700 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  605.18 699.28 605.38 700 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  607.58 699.28 607.78 700 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  257.18 699.28 257.38 700 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  609.98 699.28 610.18 700 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  612.38 699.28 612.58 700 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  614.78 699.28 614.98 700 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  254.78 699.28 254.98 700 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  617.18 699.28 617.38 700 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.58 699.28 619.78 700 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  621.98 699.28 622.18 700 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  252.38 699.28 252.58 700 ;
    END
  END instr_rdata_i[9]
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  624.38 699.28 624.58 700 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  626.78 699.28 626.98 700 ;
    END
  END instr_rvalid_i
  PIN irqs_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  629.18 699.28 629.38 700 ;
    END
  END irqs_i[0]
  PIN irqs_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  249.98 699.28 250.18 700 ;
    END
  END irqs_i[10]
  PIN irqs_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  631.58 699.28 631.78 700 ;
    END
  END irqs_i[11]
  PIN irqs_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  633.98 699.28 634.18 700 ;
    END
  END irqs_i[12]
  PIN irqs_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  636.38 699.28 636.58 700 ;
    END
  END irqs_i[13]
  PIN irqs_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  247.58 699.28 247.78 700 ;
    END
  END irqs_i[14]
  PIN irqs_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  324.38 699.28 324.58 700 ;
    END
  END irqs_i[15]
  PIN irqs_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  638.78 699.28 638.98 700 ;
    END
  END irqs_i[1]
  PIN irqs_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  641.18 699.28 641.38 700 ;
    END
  END irqs_i[2]
  PIN irqs_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  245.18 699.28 245.38 700 ;
    END
  END irqs_i[3]
  PIN irqs_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  643.58 699.28 643.78 700 ;
    END
  END irqs_i[4]
  PIN irqs_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  645.98 699.28 646.18 700 ;
    END
  END irqs_i[5]
  PIN irqs_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  648.38 699.28 648.58 700 ;
    END
  END irqs_i[6]
  PIN irqs_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  242.78 699.28 242.98 700 ;
    END
  END irqs_i[7]
  PIN irqs_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  650.78 699.28 650.98 700 ;
    END
  END irqs_i[8]
  PIN irqs_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  653.18 699.28 653.38 700 ;
    END
  END irqs_i[9]
  PIN ref_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  105.98 0 106.18 0.72 ;
    END
  END ref_clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  655.58 699.28 655.78 700 ;
    END
  END rst_ni
  PIN test_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  240.38 699.28 240.58 700 ;
    END
  END test_enable_i
  PIN timer0_irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  657.98 699.28 658.18 700 ;
    END
  END timer0_irq_i
  OBS
    LAYER Metal1 ;
     RECT  25.44 26.24 674.88 673.06 ;
    LAYER Metal2 ;
     RECT  25.34 338 25.735 338.2 ;
     RECT  25.34 357.32 25.735 360.46 ;
     RECT  25.735 269.54 25.82 277.72 ;
     RECT  25.735 307.34 25.82 315.1 ;
     RECT  25.735 338 25.82 345.76 ;
     RECT  25.735 357.32 25.82 368.44 ;
     RECT  25.735 448.46 25.82 448.66 ;
     RECT  25.735 546.32 25.82 546.52 ;
     RECT  25.82 297.68 26.215 315.1 ;
     RECT  25.735 556.82 26.215 557.02 ;
     RECT  25.735 571.94 26.215 579.7 ;
     RECT  26.215 297.68 26.3 320.14 ;
     RECT  25.82 338 26.3 348.7 ;
     RECT  25.82 357.32 26.3 376 ;
     RECT  25.735 405.62 26.3 405.82 ;
     RECT  25.735 418.22 26.3 418.42 ;
     RECT  25.82 448.46 26.3 455.8 ;
     RECT  25.735 259.46 26.515 259.66 ;
     RECT  25.735 390.5 26.515 390.7 ;
     RECT  25.735 433.34 26.515 433.54 ;
     RECT  26.3 448.46 26.515 456.22 ;
     RECT  25.735 508.94 26.515 516.7 ;
     RECT  26.215 556.82 26.515 579.7 ;
     RECT  25.735 473.66 26.655 478.9 ;
     RECT  25.82 269.54 26.695 278.56 ;
     RECT  26.3 289.7 26.695 320.14 ;
     RECT  25.82 545.48 26.695 546.52 ;
     RECT  26.3 405.62 26.78 418.42 ;
     RECT  26.78 496.76 27.175 499.06 ;
     RECT  26.515 508.1 27.175 516.7 ;
     RECT  26.695 539.18 27.175 546.52 ;
     RECT  26.3 336.74 27.205 379.78 ;
     RECT  26.695 269.54 27.26 320.14 ;
     RECT  27.205 330.02 27.26 379.78 ;
     RECT  26.78 402.68 27.26 418.42 ;
     RECT  27.175 534.14 27.26 546.52 ;
     RECT  27.26 269.54 27.685 379.78 ;
     RECT  26.515 390.5 27.685 391.54 ;
     RECT  26.655 473.66 27.74 485.83 ;
     RECT  27.175 496.76 27.74 516.7 ;
     RECT  27.26 526.16 27.74 546.52 ;
     RECT  27.74 473.66 28.095 486.04 ;
     RECT  28.095 466.73 28.135 486.04 ;
     RECT  27.74 496.76 28.135 546.52 ;
     RECT  26.515 258.62 28.22 259.66 ;
     RECT  26.515 432.5 28.22 433.54 ;
     RECT  28.22 257.36 28.7 259.66 ;
     RECT  27.685 269.54 28.7 391.54 ;
     RECT  27.26 401 28.7 421.36 ;
     RECT  28.22 432.5 28.7 436.48 ;
     RECT  26.515 447.62 28.7 456.22 ;
     RECT  28.135 466.73 28.7 546.52 ;
     RECT  28.7 256.1 29.095 391.54 ;
     RECT  28.7 466.73 29.18 547.78 ;
     RECT  26.515 556.82 29.18 580.54 ;
     RECT  28.7 400.58 29.575 421.36 ;
     RECT  28.7 432.5 29.575 456.22 ;
     RECT  29.575 400.58 29.66 456.22 ;
     RECT  29.18 466.52 29.66 547.78 ;
     RECT  29.095 251.9 29.875 391.54 ;
     RECT  29.875 251.06 30.14 391.54 ;
     RECT  29.66 400.58 30.14 547.78 ;
     RECT  29.18 556.82 30.14 584.32 ;
     RECT  30.62 110.78 31.52 110.98 ;
     RECT  30.14 251.06 32.455 584.32 ;
     RECT  31.52 110.78 33.02 111.99 ;
     RECT  32.455 251.06 33.235 587.26 ;
     RECT  33.02 110.78 33.92 118.54 ;
     RECT  34.46 130.94 35.36 131.14 ;
     RECT  33.92 110.78 35.9 119.55 ;
     RECT  35.36 129.93 35.9 131.14 ;
     RECT  39.175 599.66 39.955 599.86 ;
     RECT  39.955 598.82 40.135 599.86 ;
     RECT  35.9 110.78 40.22 131.14 ;
     RECT  33.235 251.06 40.22 588.1 ;
     RECT  40.22 251.06 41.18 588.52 ;
     RECT  40.135 598.82 41.18 607.42 ;
     RECT  41.18 251.06 42.38 607.42 ;
     RECT  42.38 247.7 43.1 607.42 ;
     RECT  40.22 107 44.06 131.14 ;
     RECT  43.1 246.86 44.54 607.42 ;
     RECT  44.06 107 45.22 131.56 ;
     RECT  45.22 107.42 45.98 131.56 ;
     RECT  44.54 244.34 46.46 607.42 ;
     RECT  45.98 107.42 46.88 133.66 ;
     RECT  46.46 239.72 47.42 607.42 ;
     RECT  47.42 236.36 49.34 607.42 ;
     RECT  49.34 235.94 50.78 607.42 ;
     RECT  50.78 235.52 51.74 607.42 ;
     RECT  46.88 107.42 52.7 134.67 ;
     RECT  51.74 235.52 54.14 610.36 ;
     RECT  52.7 107.42 56.06 139.12 ;
     RECT  54.14 235.52 57.415 612.04 ;
     RECT  57.415 235.52 58.94 614.56 ;
     RECT  59.785 210.305 60.28 210.535 ;
     RECT  56.06 106.58 60.38 139.12 ;
     RECT  60.38 106.58 61.28 141.22 ;
     RECT  61.28 106.58 62.78 142.23 ;
     RECT  62.78 106.58 63.68 156.34 ;
     RECT  58.94 232.16 63.77 614.56 ;
     RECT  63.77 232.16 63.84 614.9 ;
     RECT  63.74 168.74 64.64 168.94 ;
     RECT  63.68 106.58 65.18 157.35 ;
     RECT  65.18 103.64 65.66 157.35 ;
     RECT  64.64 167.73 65.66 168.94 ;
     RECT  65.66 103.64 66.14 168.94 ;
     RECT  63.84 232.16 66.65 614.98 ;
     RECT  66.65 231.82 66.72 614.98 ;
     RECT  66.72 231.74 69.5 614.98 ;
     RECT  60.28 209.47 69.98 210.535 ;
     RECT  69.5 231.74 71.9 617.92 ;
     RECT  66.14 102.8 73.34 168.94 ;
     RECT  69.98 209.06 73.34 210.535 ;
     RECT  73.34 102.8 75.94 169.36 ;
     RECT  75.94 103.22 77.38 169.36 ;
     RECT  71.9 231.74 79.1 622.54 ;
     RECT  79.1 231.74 81.02 625.9 ;
     RECT  77.38 103.22 81.7 164.91 ;
     RECT  81.02 231.74 81.92 632.62 ;
     RECT  85.34 648.38 86.24 649.42 ;
     RECT  81.92 231.74 86.3 633.63 ;
     RECT  81.7 103.64 86.5 164.91 ;
     RECT  73.34 209.06 86.98 211.36 ;
     RECT  86.24 648.345 87.26 649.42 ;
     RECT  86.5 106.58 87.925 164.91 ;
     RECT  86.3 231.74 88.585 635.98 ;
     RECT  87.925 106.58 90.34 163.48 ;
     RECT  88.585 227.945 90.62 635.98 ;
     RECT  87.26 647.96 90.62 649.42 ;
     RECT  90.34 148.16 91.3 163.48 ;
     RECT  90.62 647.96 91.58 651.94 ;
     RECT  91.3 148.16 92.26 152.98 ;
     RECT  91.58 647.96 92.54 655.72 ;
     RECT  92.26 152.78 93.7 152.98 ;
     RECT  86.98 209.06 94.115 210.535 ;
     RECT  90.34 106.58 94.18 138.7 ;
     RECT  90.62 227.945 94.46 637.24 ;
     RECT  94.46 227.945 94.94 638.08 ;
     RECT  92.54 647.96 94.94 656.98 ;
     RECT  94.115 209.06 95.14 210.52 ;
     RECT  94.94 227.945 95.42 656.98 ;
     RECT  95.42 223.76 99.26 656.98 ;
     RECT  99.26 223.76 102.62 659.92 ;
     RECT  102.62 222.08 103.1 659.92 ;
     RECT  94.18 107.84 103.58 138.7 ;
     RECT  103.58 107 103.78 139.12 ;
     RECT  95.14 210.32 104.06 210.52 ;
     RECT  103.1 221.24 104.06 659.92 ;
     RECT  103.78 107 110.3 131.56 ;
     RECT  110.3 104.9 110.78 131.56 ;
     RECT  104.06 210.32 112.615 659.92 ;
     RECT  110.78 104.06 113.18 131.56 ;
     RECT  112.615 210.32 113.395 662.86 ;
     RECT  113.18 104.06 114.52 133.24 ;
     RECT  113.395 210.32 116.905 663.7 ;
     RECT  116.905 202.745 117.4 663.7 ;
     RECT  117.4 201.91 117.5 663.7 ;
     RECT  117.5 198.98 118.4 663.7 ;
     RECT  118.94 144.8 119.42 148.78 ;
     RECT  119.42 141.86 119.84 148.78 ;
     RECT  118.94 186.38 119.84 186.58 ;
     RECT  119.84 186.38 119.9 187.59 ;
     RECT  118.4 197.97 119.9 663.7 ;
     RECT  119.84 141.86 120.32 149.79 ;
     RECT  114.52 103.63 121.76 133.24 ;
     RECT  120.32 141.825 121.76 149.79 ;
     RECT  121.76 103.63 121.925 149.79 ;
     RECT  119.9 186.38 123.74 663.7 ;
     RECT  121.925 103.64 124.22 149.79 ;
     RECT  123.74 184.28 125.66 663.7 ;
     RECT  125.66 179.66 127.1 663.7 ;
     RECT  127.1 177.98 127.58 663.7 ;
     RECT  127.58 177.98 128.06 664.54 ;
     RECT  124.22 103.64 129.02 152.98 ;
     RECT  129.02 103.64 133.82 160.96 ;
     RECT  133.82 103.64 135.145 168.94 ;
     RECT  128.06 177.98 135.145 672.1 ;
     RECT  135.145 103.64 135.94 672.1 ;
     RECT  135.94 104.06 138.34 672.1 ;
     RECT  138.34 106.58 144.58 672.1 ;
     RECT  144.58 106.58 151.1 671.68 ;
     RECT  151.1 103.22 158.78 671.68 ;
     RECT  158.78 99.86 160.42 671.68 ;
     RECT  160.42 99.86 166.18 671.26 ;
     RECT  166.18 100.28 167.62 671.26 ;
     RECT  167.62 100.7 176 671.26 ;
     RECT  176 100.7 177.5 671.43 ;
     RECT  177.5 100.28 179.42 671.43 ;
     RECT  179.42 99.86 183.445 671.43 ;
     RECT  183.445 99.86 192.595 670.42 ;
     RECT  192.595 99.86 201.45 671.26 ;
     RECT  201.45 99.86 210.62 670.84 ;
     RECT  210.62 99.86 213.98 672.52 ;
     RECT  213.98 99.44 220.9 672.52 ;
     RECT  220.9 99.86 222.34 672.52 ;
     RECT  222.34 100.7 223.3 672.52 ;
     RECT  221.18 697.52 223.58 697.72 ;
     RECT  223.3 130.52 225.98 672.52 ;
     RECT  223.3 100.7 228.565 119.55 ;
     RECT  228.565 100.7 230.02 118.12 ;
     RECT  230.02 107.42 231.94 118.12 ;
     RECT  225.98 130.52 236.06 680.5 ;
     RECT  236.06 126.74 240.58 680.5 ;
     RECT  240.58 130.94 241.06 680.5 ;
     RECT  241.06 131.36 247.3 680.5 ;
     RECT  223.58 696.68 250.46 697.72 ;
     RECT  247.3 131.36 251.14 142.9 ;
     RECT  247.3 152.61 254.02 680.5 ;
     RECT  254.02 152.61 254.485 214.72 ;
     RECT  254.485 153.2 254.98 214.72 ;
     RECT  251.14 137.225 255.875 142.9 ;
     RECT  255.875 138.06 256.325 142.9 ;
     RECT  254.98 153.62 256.42 214.72 ;
     RECT  231.94 107.42 256.9 107.62 ;
     RECT  256.325 138.08 256.9 142.9 ;
     RECT  256.9 142.7 257.38 142.9 ;
     RECT  254.02 225.02 257.845 680.5 ;
     RECT  256.42 153.62 257.86 154.24 ;
     RECT  250.46 694.16 259.58 697.72 ;
     RECT  257.845 228.38 261.22 680.5 ;
     RECT  256.42 167.73 266.3 214.72 ;
     RECT  261.22 228.38 266.3 328.12 ;
     RECT  266.3 136.36 268.7 136.56 ;
     RECT  266.3 147.7 268.7 149.58 ;
     RECT  266.3 159.04 268.7 328.12 ;
     RECT  268.7 131.32 269.675 138.66 ;
     RECT  268.7 147.7 269.675 328.12 ;
     RECT  261.22 336.7 269.675 680.5 ;
     RECT  269.675 131.32 271.675 680.5 ;
     RECT  271.675 131.31 273.98 680.5 ;
     RECT  271.1 113.68 275.9 113.88 ;
     RECT  259.58 694.16 276.58 698.98 ;
     RECT  275.9 109.9 277.34 113.88 ;
     RECT  273.98 122.92 277.34 680.5 ;
     RECT  277.34 109.9 279.275 680.5 ;
     RECT  279.275 109.06 282.34 680.5 ;
     RECT  282.34 109.06 282.495 409.56 ;
     RECT  282.495 105.28 283.1 409.56 ;
     RECT  282.34 421.58 293.18 680.5 ;
     RECT  283.1 100.66 298.46 409.56 ;
     RECT  298.46 97.72 301.82 409.56 ;
     RECT  293.18 421.58 301.82 687.64 ;
     RECT  301.82 97.72 306.14 687.64 ;
     RECT  306.14 96.46 307.78 687.64 ;
     RECT  307.78 96.46 310.18 426.36 ;
     RECT  310.18 96.88 317.38 426.36 ;
     RECT  307.78 435.44 317.86 687.64 ;
     RECT  317.38 97.72 318.45 426.36 ;
     RECT  318.45 98.56 326.02 426.36 ;
     RECT  326.02 100.24 330.82 426.36 ;
     RECT  330.82 101.465 331.36 426.36 ;
     RECT  331.36 101.5 341.18 426.36 ;
     RECT  341.18 101.5 341.66 426.78 ;
     RECT  341.66 101.08 347.42 426.78 ;
     RECT  347.42 98.56 350.795 426.78 ;
     RECT  350.795 97.13 360.86 426.78 ;
     RECT  360.86 93.94 361.82 426.78 ;
     RECT  361.82 93.52 363.74 426.78 ;
     RECT  363.74 93.1 366.62 426.78 ;
     RECT  366.62 93.1 373.54 427.2 ;
     RECT  373.54 93.52 375.46 427.2 ;
     RECT  375.46 96.46 389.66 427.2 ;
     RECT  317.86 440.06 394.18 687.64 ;
     RECT  389.66 96.46 395.14 429.3 ;
     RECT  276.58 696.68 403.58 698.98 ;
     RECT  395.14 97.72 404.06 429.3 ;
     RECT  404.06 97.3 405.5 429.3 ;
     RECT  405.5 97.3 417.02 430.56 ;
     RECT  417.02 96.88 419.42 430.56 ;
     RECT  394.18 440.06 419.42 680.5 ;
     RECT  419.42 96.88 421.54 680.5 ;
     RECT  421.54 97.72 423.46 680.5 ;
     RECT  403.58 691.22 432.1 698.98 ;
     RECT  432.1 691.22 434.02 698.56 ;
     RECT  423.46 100.66 446.3 680.5 ;
     RECT  434.02 691.22 448.9 691.42 ;
     RECT  446.3 97.3 453.22 680.5 ;
     RECT  453.22 98.14 455.14 680.5 ;
     RECT  455.14 100.66 461.86 680.5 ;
     RECT  461.86 103.6 465.98 680.5 ;
     RECT  456.38 692.06 465.98 692.26 ;
     RECT  465.98 103.6 472.42 692.26 ;
     RECT  472.42 105.28 473.86 675.46 ;
     RECT  473.86 106.54 481.54 675.46 ;
     RECT  472.42 684.08 482.5 692.26 ;
     RECT  482.5 692.06 486.82 692.26 ;
     RECT  481.54 106.54 488.74 426.36 ;
     RECT  481.54 439.6 494.5 675.46 ;
     RECT  488.74 107.8 501.98 426.36 ;
     RECT  494.5 440.02 504.38 675.46 ;
     RECT  501.98 104.86 506.795 426.36 ;
     RECT  506.795 104.69 514.24 426.36 ;
     RECT  514.24 105.7 514.46 426.36 ;
     RECT  514.46 105.7 515.62 426.78 ;
     RECT  504.38 435.82 518.98 675.46 ;
     RECT  518.98 435.82 525.5 674.2 ;
     RECT  515.62 107.38 525.98 426.78 ;
     RECT  525.98 104.86 531.275 426.78 ;
     RECT  525.5 435.4 533.38 674.2 ;
     RECT  531.275 104.69 540.86 426.78 ;
     RECT  540.86 102.34 544.235 426.78 ;
     RECT  533.38 440.02 545.66 674.2 ;
     RECT  544.235 101.5 551.39 426.78 ;
     RECT  551.39 101.465 551.68 426.78 ;
     RECT  551.68 102.34 555.46 426.78 ;
     RECT  555.46 104.02 556.42 425.52 ;
     RECT  556.42 104.02 557.38 425.1 ;
     RECT  557.38 105.28 560.26 425.1 ;
     RECT  560.26 105.28 566.795 424.68 ;
     RECT  545.66 440.02 566.98 675.04 ;
     RECT  566.98 440.02 572.26 674.62 ;
     RECT  572.26 440.02 572.74 674.2 ;
     RECT  566.795 104.69 574.24 424.68 ;
     RECT  574.24 108.22 585.22 424.68 ;
     RECT  585.22 108.22 585.7 424.26 ;
     RECT  572.74 440.02 586.66 672.52 ;
     RECT  585.7 108.64 587.14 424.26 ;
     RECT  587.14 109.48 589.06 424.26 ;
     RECT  585.98 691.22 590.78 691.42 ;
     RECT  590.78 691.22 593.18 693.94 ;
     RECT  586.66 440.86 597.94 672.52 ;
     RECT  597.94 514.82 600.58 672.52 ;
     RECT  589.06 112.25 600.64 424.26 ;
     RECT  600.64 113.26 601.54 424.26 ;
     RECT  601.54 114.94 602.98 424.26 ;
     RECT  593.18 691.22 602.98 695.2 ;
     RECT  597.94 440.86 604.9 504.52 ;
     RECT  600.58 514.82 604.9 670.84 ;
     RECT  602.98 114.94 606.34 421.74 ;
     RECT  604.9 451.82 606.82 496.54 ;
     RECT  606.82 451.82 607.3 496.12 ;
     RECT  607.3 455.6 607.78 496.12 ;
     RECT  607.78 456.44 608.26 496.12 ;
     RECT  608.26 456.44 609.7 495.7 ;
     RECT  606.34 114.94 610.18 417.96 ;
     RECT  602.98 693.32 611.42 695.2 ;
     RECT  609.7 457.28 611.62 495.7 ;
     RECT  611.62 457.28 612.1 494.44 ;
     RECT  612.1 461.9 612.34 494.44 ;
     RECT  612.34 462.74 612.82 494.44 ;
     RECT  612.82 462.74 613.06 489.4 ;
     RECT  613.06 464 613.54 489.4 ;
     RECT  613.54 464 613.78 488.56 ;
     RECT  604.9 440.86 614.02 441.06 ;
     RECT  613.78 471.14 614.5 488.56 ;
     RECT  611.42 692.9 614.78 695.2 ;
     RECT  614.5 471.14 614.98 486.04 ;
     RECT  604.9 515.49 616.405 670.84 ;
     RECT  614.98 471.56 616.42 486.04 ;
     RECT  616.42 473.66 617.38 486.04 ;
     RECT  617.38 473.66 617.86 485.2 ;
     RECT  617.86 482.06 618.82 485.2 ;
     RECT  618.82 483.74 619.3 485.2 ;
     RECT  619.3 485 619.54 485.2 ;
     RECT  616.405 516.92 619.78 670.84 ;
     RECT  614.78 692.48 620.26 695.2 ;
     RECT  610.18 114.94 621.22 417.12 ;
     RECT  621.22 416.92 621.7 417.12 ;
     RECT  620.26 692.9 622.66 695.2 ;
     RECT  621.22 114.94 624.86 403.68 ;
     RECT  619.78 518.6 625.06 670.84 ;
     RECT  622.66 692.9 626.02 693.52 ;
     RECT  624.86 113.68 626.78 403.68 ;
     RECT  626.02 692.9 626.98 693.1 ;
     RECT  625.06 519.86 627.94 670.84 ;
     RECT  626.78 112.42 628.235 403.68 ;
     RECT  627.94 519.86 631.285 663.7 ;
     RECT  631.285 520.7 634.66 663.7 ;
     RECT  628.235 112.25 635.68 403.68 ;
     RECT  635.68 113.26 637.06 403.68 ;
     RECT  634.66 521.12 638.02 663.7 ;
     RECT  638.02 524.48 638.5 663.7 ;
     RECT  638.5 530.61 638.98 663.7 ;
     RECT  638.98 530.61 642.805 662.86 ;
     RECT  637.06 116.2 642.82 403.68 ;
     RECT  642.805 531.62 645.22 662.86 ;
     RECT  642.82 120.4 647.62 403.68 ;
     RECT  647.62 127.37 649.06 403.68 ;
     RECT  649.06 127.37 649.54 388.98 ;
     RECT  649.54 127.37 650.02 386.04 ;
     RECT  650.02 138.46 650.5 386.04 ;
     RECT  650.5 138.46 650.98 143.7 ;
     RECT  650.5 154 650.98 386.04 ;
     RECT  650.02 127.37 651.04 128.58 ;
     RECT  651.04 128.38 651.94 128.58 ;
     RECT  645.22 531.62 652.105 659.92 ;
     RECT  650.98 138.46 652.48 139.67 ;
     RECT  650.98 154 652.9 385.2 ;
     RECT  652.48 138.46 653.38 138.66 ;
     RECT  652.105 530.345 656.26 659.92 ;
     RECT  656.26 542.12 656.74 659.92 ;
     RECT  656.74 659.72 658.66 659.92 ;
     RECT  652.9 154 659.14 381 ;
     RECT  656.26 530.345 659.555 531.82 ;
     RECT  659.14 154 659.62 154.2 ;
     RECT  659.555 531.18 660.005 531.82 ;
     RECT  659.14 162.82 660.58 381 ;
     RECT  660.005 531.2 660.58 531.82 ;
     RECT  656.74 542.12 660.58 646.9 ;
     RECT  660.58 162.82 661.06 230.39 ;
     RECT  661.06 162.82 661.54 172.26 ;
     RECT  660.58 542.12 661.54 643.54 ;
     RECT  661.54 166.6 662.02 172.26 ;
     RECT  661.06 181.3 662.02 230.39 ;
     RECT  660.58 240.77 662.02 381 ;
     RECT  662.02 191.38 662.5 206.7 ;
     RECT  662.02 240.77 662.5 336.48 ;
     RECT  662.02 358.96 662.5 381 ;
     RECT  661.54 542.12 662.5 635.98 ;
     RECT  662.02 218.09 662.56 230.39 ;
     RECT  662.5 252.665 662.98 336.48 ;
     RECT  662.5 542.12 662.98 619.18 ;
     RECT  662.02 169.505 663.04 172.26 ;
     RECT  662.5 191.38 663.46 200.82 ;
     RECT  662.98 309.4 663.46 336.48 ;
     RECT  662.56 222.04 663.52 230.39 ;
     RECT  662.5 240.77 663.52 241.98 ;
     RECT  662.98 252.665 663.52 290.7 ;
     RECT  662.5 361.73 663.52 377.22 ;
     RECT  663.04 169.54 663.94 172.26 ;
     RECT  662.5 630.32 663.94 635.98 ;
     RECT  663.46 191.38 664 192.59 ;
     RECT  663.52 255.22 664 290.7 ;
     RECT  663.46 324.1 664 336.48 ;
     RECT  663.52 222.04 664.42 229.38 ;
     RECT  663.52 241.78 664.42 241.98 ;
     RECT  664 255.22 664.42 262.98 ;
     RECT  664 287.14 664.42 290.7 ;
     RECT  664 324.1 664.42 324.72 ;
     RECT  663.52 368.62 664.42 377.22 ;
     RECT  663.94 630.32 664.42 630.52 ;
     RECT  664 191.38 664.9 191.58 ;
     RECT  664.42 262.78 664.9 262.98 ;
     RECT  664 277.9 664.9 278.1 ;
     RECT  664.42 290.5 664.9 290.7 ;
     RECT  664 336.28 664.9 336.48 ;
     RECT  662.98 543.38 666.34 619.18 ;
     RECT  666.34 545.06 670.18 619.18 ;
     RECT  670.18 548.84 671.125 619.18 ;
     RECT  671.125 569.84 671.62 619.18 ;
     RECT  671.62 569.84 672.1 609.52 ;
     RECT  671.125 548.84 673.54 560.38 ;
     RECT  673.54 555.98 674.5 560.38 ;
     RECT  672.1 569.84 674.5 579.28 ;
     RECT  672.1 588.74 674.5 609.52 ;
    LAYER Metal3 ;
     RECT  22.46 0.32 24.1 0.42 ;
     RECT  101.66 0.32 103.3 0.42 ;
     RECT  21.98 0.42 24.58 0.94 ;
     RECT  101.18 0.42 103.78 0.94 ;
     RECT  370.94 93.1 371.14 93.52 ;
     RECT  361.82 93.52 371.14 93.94 ;
     RECT  360.86 93.94 374.5 96.16 ;
     RECT  360.86 96.16 374.98 96.46 ;
     RECT  309.98 96.46 310.18 96.88 ;
     RECT  360.86 96.46 389.86 96.88 ;
     RECT  309.02 96.88 312.1 97.3 ;
     RECT  360.86 96.88 394.66 97.3 ;
     RECT  309.02 97.3 315.46 97.72 ;
     RECT  357.98 97.3 394.66 97.72 ;
     RECT  417.02 96.88 421.54 97.72 ;
     RECT  446.3 97.3 446.5 97.72 ;
     RECT  357.5 97.72 394.66 98.14 ;
     RECT  446.3 97.72 450.82 98.14 ;
     RECT  309.02 97.72 317.86 98.56 ;
     RECT  354.14 98.14 397.06 98.56 ;
     RECT  197.66 99.44 197.86 99.86 ;
     RECT  213.98 99.44 218.5 99.86 ;
     RECT  309.02 98.56 326.02 100.24 ;
     RECT  162.14 99.44 169.54 100.28 ;
     RECT  182.78 99.44 182.98 100.28 ;
     RECT  197.66 99.86 202.18 100.28 ;
     RECT  213.98 99.86 222.34 100.28 ;
     RECT  417.02 97.72 424.42 100.66 ;
     RECT  446.3 98.14 452.26 100.66 ;
     RECT  213.5 100.28 222.34 100.7 ;
     RECT  283.1 100.66 283.3 101.08 ;
     RECT  298.46 97.72 298.66 101.08 ;
     RECT  349.82 98.56 397.54 101.08 ;
     RECT  417.02 100.66 452.26 101.08 ;
     RECT  309.02 100.24 330.82 101.5 ;
     RECT  341.66 101.08 397.54 101.5 ;
     RECT  407.42 101.08 452.26 101.5 ;
     RECT  550.46 101.08 550.66 101.5 ;
     RECT  407.42 101.5 452.74 102.34 ;
     RECT  213.5 100.7 230.02 103 ;
     RECT  67.1 103.22 67.3 103.64 ;
     RECT  80.06 103.22 83.62 103.64 ;
     RECT  158.78 100.28 202.66 103.64 ;
     RECT  213.5 103 225.7 103.64 ;
     RECT  544.22 101.5 552.58 104.44 ;
     RECT  127.58 103.64 136.42 104.48 ;
     RECT  283.1 101.08 298.66 104.86 ;
     RECT  309.02 101.5 397.54 104.86 ;
     RECT  407.42 102.34 455.62 104.86 ;
     RECT  544.22 104.44 557.38 104.86 ;
     RECT  105.02 102.8 105.22 104.9 ;
     RECT  283.1 104.86 461.38 105.28 ;
     RECT  501.98 104.86 502.18 105.28 ;
     RECT  525.98 104.86 526.18 105.28 ;
     RECT  540.86 104.86 557.38 105.28 ;
     RECT  573.98 104.86 574.18 105.28 ;
     RECT  472.22 103.6 472.42 105.7 ;
     RECT  525.98 105.28 574.18 105.7 ;
     RECT  282.62 105.28 461.38 106.12 ;
     RECT  471.74 105.7 472.42 106.12 ;
     RECT  501.98 105.28 508.42 106.12 ;
     RECT  127.58 104.48 136.9 106.58 ;
     RECT  127.58 106.58 143.14 107 ;
     RECT  153.02 103.64 225.7 107 ;
     RECT  501.98 106.12 509.38 107.38 ;
     RECT  525.98 105.7 575.14 107.38 ;
     RECT  65.18 103.64 83.62 107.42 ;
     RECT  105.02 104.9 110.5 107.42 ;
     RECT  282.62 106.12 472.42 107.8 ;
     RECT  488.54 106.54 488.74 107.8 ;
     RECT  40.22 107 40.42 107.84 ;
     RECT  53.66 107 53.86 107.84 ;
     RECT  63.74 107.42 83.62 107.84 ;
     RECT  105.02 107.42 112.9 107.84 ;
     RECT  501.98 107.38 575.14 108.22 ;
     RECT  40.22 107.84 41.38 108.26 ;
     RECT  53.66 107.84 84.1 108.26 ;
     RECT  98.78 107.84 112.9 108.26 ;
     RECT  282.62 107.8 488.74 108.64 ;
     RECT  501.98 108.22 578.98 108.64 ;
     RECT  282.62 108.64 587.14 109.48 ;
     RECT  282.62 109.48 589.06 109.9 ;
     RECT  40.22 108.26 84.1 110.78 ;
     RECT  98.3 108.26 112.9 110.78 ;
     RECT  127.58 107 225.7 110.98 ;
     RECT  40.22 110.78 112.9 111.2 ;
     RECT  281.66 109.9 589.06 112.42 ;
     RECT  34.94 111.2 112.9 112.46 ;
     RECT  127.58 110.98 223.3 112.46 ;
     RECT  281.66 112.42 592.9 112.84 ;
     RECT  626.78 112.42 626.98 112.84 ;
     RECT  626.78 112.84 633.22 113.26 ;
     RECT  281.66 112.84 599.62 115.36 ;
     RECT  626.78 113.26 637.06 115.78 ;
     RECT  626.78 115.78 637.54 116.2 ;
     RECT  271.1 113.68 271.3 116.62 ;
     RECT  281.66 115.36 602.98 116.62 ;
     RECT  271.1 116.62 604.42 117.46 ;
     RECT  617.66 116.2 642.82 117.46 ;
     RECT  34.94 112.46 223.3 118.96 ;
     RECT  271.1 117.46 642.82 120.4 ;
     RECT  35.9 118.96 223.3 121.9 ;
     RECT  35.9 121.9 183.46 124 ;
     RECT  271.1 120.4 647.62 127.96 ;
     RECT  236.54 126.74 236.74 129.68 ;
     RECT  193.34 121.9 223.3 130.52 ;
     RECT  236.54 129.68 240.1 130.52 ;
     RECT  35.9 124 182.5 130.72 ;
     RECT  193.34 130.52 240.1 130.94 ;
     RECT  271.1 127.96 650.02 131.1 ;
     RECT  35.9 130.72 61.06 131.14 ;
     RECT  271.1 131.1 649.06 131.32 ;
     RECT  193.34 130.94 241.06 131.36 ;
     RECT  256.7 107.42 256.9 131.36 ;
     RECT  44.06 131.14 61.06 131.56 ;
     RECT  71.42 130.72 182.5 131.56 ;
     RECT  71.42 131.56 96.1 133.24 ;
     RECT  113.18 131.56 182.5 133.24 ;
     RECT  120.86 133.24 182.5 133.66 ;
     RECT  50.3 131.56 61.06 134.08 ;
     RECT  121.34 133.66 182.5 134.3 ;
     RECT  193.34 131.36 256.9 134.3 ;
     RECT  71.42 133.24 94.66 137.86 ;
     RECT  71.42 137.86 94.18 138.28 ;
     RECT  121.34 134.3 256.9 138.28 ;
     RECT  53.66 134.08 61.06 139.12 ;
     RECT  71.42 138.28 93.7 139.12 ;
     RECT  71.42 139.12 82.66 141.44 ;
     RECT  268.7 131.32 649.06 146.02 ;
     RECT  121.34 138.28 254.02 149.2 ;
     RECT  65.18 141.44 82.66 149.62 ;
     RECT  127.1 149.2 254.02 152.14 ;
     RECT  93.5 139.12 93.7 152.98 ;
     RECT  81.98 149.62 82.66 153.2 ;
     RECT  128.06 152.14 254.02 153.2 ;
     RECT  268.7 146.02 650.5 153.58 ;
     RECT  268.7 153.58 657.7 154 ;
     RECT  668.54 31.46 668.74 154 ;
     RECT  128.06 153.2 254.98 154.24 ;
     RECT  81.98 153.2 87.46 155.92 ;
     RECT  268.7 154 668.74 156.3 ;
     RECT  65.18 149.62 72.1 159.92 ;
     RECT  81.98 155.92 85.54 159.92 ;
     RECT  129.5 154.24 254.98 160.34 ;
     RECT  65.18 159.92 85.54 160.54 ;
     RECT  129.5 160.34 256.42 160.96 ;
     RECT  65.18 160.54 82.18 164.74 ;
     RECT  272.54 156.3 668.74 165.96 ;
     RECT  65.18 164.74 73.54 168.52 ;
     RECT  274.46 165.96 668.74 168.9 ;
     RECT  65.66 168.52 73.54 168.94 ;
     RECT  73.34 168.94 73.54 169.36 ;
     RECT  129.98 160.96 256.42 173.78 ;
     RECT  129.98 173.78 256.9 178.82 ;
     RECT  129.98 178.82 257.38 179.24 ;
     RECT  274.94 168.9 668.74 184.66 ;
     RECT  129.5 179.24 257.38 187.22 ;
     RECT  127.1 187.22 257.38 188.06 ;
     RECT  127.1 188.06 262.66 193.06 ;
     RECT  273.02 184.66 668.74 193.06 ;
     RECT  127.1 193.06 668.74 194.36 ;
     RECT  121.82 194.36 668.74 198.56 ;
     RECT  94.94 209.48 95.14 211.16 ;
     RECT  119.42 198.56 668.74 214.52 ;
     RECT  107.42 214.1 107.62 216.2 ;
     RECT  107.42 216.2 108.1 220.82 ;
     RECT  118.94 214.52 668.74 220.82 ;
     RECT  86.78 211.16 95.14 221.24 ;
     RECT  107.42 220.82 668.74 221.24 ;
     RECT  69.98 231.74 70.18 232.16 ;
     RECT  46.46 219.56 46.66 235.52 ;
     RECT  58.94 232.16 59.14 235.52 ;
     RECT  69.98 232.16 74.5 236.36 ;
     RECT  86.78 221.24 668.74 236.36 ;
     RECT  46.46 235.52 59.14 236.78 ;
     RECT  69.98 236.36 668.74 236.78 ;
     RECT  46.46 236.78 668.74 244.34 ;
     RECT  44.54 244.34 668.74 246.86 ;
     RECT  32.06 251.48 32.26 254 ;
     RECT  43.1 246.86 668.74 254 ;
     RECT  32.06 254 668.74 254.84 ;
     RECT  28.22 254.84 668.74 266.8 ;
     RECT  29.66 266.8 668.74 271 ;
     RECT  30.62 271 668.74 314.9 ;
     RECT  27.74 314.9 668.74 319.94 ;
     RECT  26.3 319.94 668.74 338 ;
     RECT  25.34 338 668.74 360.46 ;
     RECT  29.66 360.46 668.74 381.84 ;
     RECT  29.66 381.84 650.98 383.36 ;
     RECT  28.7 383.36 650.98 385.2 ;
     RECT  28.7 385.2 649.06 388.4 ;
     RECT  28.22 388.4 649.06 390.7 ;
     RECT  29.66 390.7 649.06 399.9 ;
     RECT  29.66 399.9 627.46 400.58 ;
     RECT  28.7 400.58 627.46 400.74 ;
     RECT  644.06 399.9 649.06 400.74 ;
     RECT  28.7 400.74 624.1 402 ;
     RECT  28.7 402 621.7 403.26 ;
     RECT  648.86 400.74 649.06 403.68 ;
     RECT  28.7 403.26 588.58 404.52 ;
     RECT  598.46 403.26 621.7 404.52 ;
     RECT  28.7 404.52 566.5 404.94 ;
     RECT  581.18 404.52 586.66 405.36 ;
     RECT  28.7 404.94 560.26 406.04 ;
     RECT  25.82 406.04 560.26 409.56 ;
     RECT  25.82 409.56 282.34 410.44 ;
     RECT  292.22 409.56 560.26 411.24 ;
     RECT  292.22 411.24 318.82 411.66 ;
     RECT  331.58 411.24 560.26 414.18 ;
     RECT  331.58 414.18 348.58 414.6 ;
     RECT  358.94 414.18 560.26 415.02 ;
     RECT  602.78 404.52 621.7 417.12 ;
     RECT  331.58 414.6 347.62 417.54 ;
     RECT  292.22 411.66 316.42 417.7 ;
     RECT  359.42 415.02 560.26 418.38 ;
     RECT  336.38 417.54 347.62 420.06 ;
     RECT  29.66 410.44 282.34 420.1 ;
     RECT  359.42 418.38 546.34 421.74 ;
     RECT  602.78 417.12 614.02 421.74 ;
     RECT  366.62 421.74 546.34 423.84 ;
     RECT  602.78 421.74 602.98 424.26 ;
     RECT  585.02 405.36 586.66 424.68 ;
     RECT  341.18 420.06 347.62 425.1 ;
     RECT  556.22 418.38 560.26 425.1 ;
     RECT  341.18 425.1 343.78 425.52 ;
     RECT  556.22 425.1 556.42 425.52 ;
     RECT  341.18 425.52 341.38 426.78 ;
     RECT  366.62 423.84 366.82 427.2 ;
     RECT  30.14 420.1 282.34 429.14 ;
     RECT  292.7 417.7 316.42 429.14 ;
     RECT  30.14 429.14 316.42 435.44 ;
     RECT  30.14 435.44 317.86 436.28 ;
     RECT  383.42 423.84 546.34 436.7 ;
     RECT  28.7 436.28 317.86 439.42 ;
     RECT  613.82 421.74 614.02 441.06 ;
     RECT  380.06 436.7 546.34 441.32 ;
     RECT  336.38 441.32 336.58 441.74 ;
     RECT  380.06 441.32 550.66 442.16 ;
     RECT  29.18 439.42 317.86 443.42 ;
     RECT  565.34 442.58 565.54 443.42 ;
     RECT  586.46 424.68 586.66 443.42 ;
     RECT  336.38 441.74 344.74 443.84 ;
     RECT  363.26 443.42 363.46 443.84 ;
     RECT  374.3 442.16 550.66 443.84 ;
     RECT  563.9 443.42 565.54 443.84 ;
     RECT  579.26 443.42 586.66 443.84 ;
     RECT  363.26 443.84 591.46 444.26 ;
     RECT  363.26 444.26 596.74 445.1 ;
     RECT  29.18 443.42 323.62 446.36 ;
     RECT  333.98 443.84 351.46 446.36 ;
     RECT  29.18 446.36 351.46 448.04 ;
     RECT  362.3 445.1 596.74 448.04 ;
     RECT  29.18 448.04 596.74 448.46 ;
     RECT  29.18 448.46 597.22 448.88 ;
     RECT  29.18 448.88 604.9 451.82 ;
     RECT  29.18 451.82 607.3 453.92 ;
     RECT  26.78 453.92 607.3 455.8 ;
     RECT  29.18 455.8 607.3 456.44 ;
     RECT  29.18 456.44 609.7 457.28 ;
     RECT  29.18 457.28 612.1 466.94 ;
     RECT  29.18 466.94 613.06 467.36 ;
     RECT  29.18 467.36 613.54 474.5 ;
     RECT  28.7 474.5 613.54 478.06 ;
     RECT  29.18 478.06 613.54 482.06 ;
     RECT  29.18 482.06 618.82 486.04 ;
     RECT  29.18 486.04 612.1 493.6 ;
     RECT  638.3 491.72 638.5 494.24 ;
     RECT  29.18 493.6 611.62 495.7 ;
     RECT  29.18 495.7 607.3 496.12 ;
     RECT  29.18 496.12 604.9 496.34 ;
     RECT  28.7 496.34 604.9 497.8 ;
     RECT  29.18 497.8 604.9 501.58 ;
     RECT  29.66 501.58 604.9 504.52 ;
     RECT  631.1 494.24 638.5 515.24 ;
     RECT  29.66 504.52 601.06 515.66 ;
     RECT  29.66 515.66 609.22 516.08 ;
     RECT  29.66 516.08 610.18 516.5 ;
     RECT  28.7 516.5 610.18 516.92 ;
     RECT  631.1 515.24 641.86 517.76 ;
     RECT  627.26 517.76 641.86 518.3 ;
     RECT  28.7 516.92 614.02 519.44 ;
     RECT  627.26 518.3 642.34 519.44 ;
     RECT  28.7 519.44 642.34 523.64 ;
     RECT  27.74 523.64 642.34 528.26 ;
     RECT  27.26 528.26 642.34 529.1 ;
     RECT  27.26 529.1 643.3 531.4 ;
     RECT  30.14 531.4 643.3 531.62 ;
     RECT  30.14 531.62 645.7 532.04 ;
     RECT  30.14 532.04 652.42 534.34 ;
     RECT  31.58 534.34 652.42 534.56 ;
     RECT  31.58 534.56 653.86 535.4 ;
     RECT  31.58 535.4 655.78 541.7 ;
     RECT  668.54 381.84 668.74 541.7 ;
     RECT  31.58 541.7 668.74 547.58 ;
     RECT  28.7 547.58 668.74 554.08 ;
     RECT  29.66 554.08 668.74 568.7 ;
     RECT  29.18 568.7 668.74 584.32 ;
     RECT  40.22 584.32 668.74 588.52 ;
     RECT  43.1 588.52 668.74 591.88 ;
     RECT  45.02 591.88 668.74 592.52 ;
     RECT  45.02 592.52 670.18 595.24 ;
     RECT  45.02 595.24 668.74 603.86 ;
     RECT  43.1 603.86 668.74 607.42 ;
     RECT  51.74 607.42 668.74 609.32 ;
     RECT  51.74 609.32 669.22 610.36 ;
     RECT  57.5 610.36 669.22 613.72 ;
     RECT  71.9 613.72 669.22 614.14 ;
     RECT  57.5 613.72 57.7 614.56 ;
     RECT  71.9 614.14 668.74 622.54 ;
     RECT  79.1 622.54 668.74 625.9 ;
     RECT  82.46 625.9 668.74 633.04 ;
     RECT  86.3 633.04 668.74 635.98 ;
     RECT  92.54 635.98 668.74 648.38 ;
     RECT  91.58 648.38 668.74 654.88 ;
     RECT  95.42 654.88 99.46 655.72 ;
     RECT  109.82 654.88 668.74 659.5 ;
     RECT  99.26 655.72 99.46 659.92 ;
     RECT  113.18 659.5 668.74 659.92 ;
     RECT  114.14 659.92 668.74 662.44 ;
     RECT  114.14 662.44 115.3 662.86 ;
     RECT  125.66 662.44 668.74 663.28 ;
     RECT  114.62 662.86 115.3 663.7 ;
     RECT  129.5 663.28 668.74 663.7 ;
     RECT  129.98 663.7 668.74 666.22 ;
     RECT  129.98 666.22 164.26 667.48 ;
     RECT  174.62 666.22 668.74 667.9 ;
     RECT  174.62 667.9 194.5 668.32 ;
     RECT  129.98 667.48 159.94 669.58 ;
     RECT  175.1 668.32 194.5 670 ;
     RECT  175.1 670 175.3 670.42 ;
     RECT  188.54 670 194.5 670.42 ;
     RECT  204.38 667.9 668.74 670.42 ;
     RECT  129.98 669.58 130.66 670.84 ;
     RECT  141.02 669.58 159.94 670.84 ;
     RECT  221.18 670.42 668.74 670.84 ;
     RECT  130.46 670.84 130.66 671.26 ;
     RECT  151.1 670.84 158.02 671.26 ;
     RECT  194.3 670.42 194.5 671.26 ;
     RECT  221.18 670.84 264.58 671.26 ;
     RECT  284.06 670.84 320.74 671.26 ;
     RECT  151.1 671.26 151.3 671.68 ;
     RECT  359.9 670.84 526.18 672.1 ;
     RECT  210.62 670.42 210.82 672.52 ;
     RECT  536.54 670.84 668.74 673.78 ;
     RECT  367.58 672.1 526.18 674.2 ;
     RECT  392.54 674.2 526.18 675.04 ;
     RECT  545.66 673.78 668.74 675.04 ;
     RECT  507.26 675.04 526.18 681.14 ;
     RECT  392.54 675.04 448.9 684.5 ;
     RECT  290.78 671.26 320.74 687.44 ;
     RECT  331.58 670.84 346.18 687.44 ;
     RECT  549.98 675.04 668.74 687.64 ;
     RECT  507.26 681.14 533.38 688.7 ;
     RECT  367.58 674.2 374.5 691.22 ;
     RECT  391.1 684.5 448.9 691.22 ;
     RECT  458.78 675.04 495.94 691.22 ;
     RECT  507.26 688.7 535.78 691.22 ;
     RECT  290.78 687.44 346.18 691.64 ;
     RECT  225.98 671.26 264.58 693.32 ;
     RECT  225.98 693.32 271.78 694.16 ;
     RECT  225.98 694.16 276.58 694.58 ;
     RECT  290.78 691.64 350.98 695 ;
     RECT  367.58 691.22 535.78 695 ;
     RECT  290.78 695 535.78 695.42 ;
     RECT  549.98 687.64 660.58 695.42 ;
     RECT  225.98 694.58 278.98 695.84 ;
     RECT  290.78 695.42 660.58 695.84 ;
     RECT  225.98 695.84 660.58 696.68 ;
     RECT  223.58 696.68 660.58 697.52 ;
     RECT  221.18 697.52 660.58 697.94 ;
     RECT  218.78 697.94 660.58 699.3 ;
     RECT  226.46 699.3 228.1 699.4 ;
     RECT  246.14 699.3 259.3 699.4 ;
     RECT  303.26 699.3 312.1 699.4 ;
     RECT  339.26 699.3 340.9 699.4 ;
     RECT  389.66 699.3 398.5 699.4 ;
     RECT  411.26 699.3 441.22 699.4 ;
     RECT  461.66 699.3 465.7 699.4 ;
     RECT  476.06 699.3 494.5 699.4 ;
     RECT  507.26 699.3 520.42 699.4 ;
     RECT  584.06 699.3 642.34 699.4 ;
    LAYER Metal4 ;
     RECT  25.82 406.04 28.7 406.24 ;
     RECT  28.22 527 28.7 527.2 ;
     RECT  30.14 468.2 30.62 468.4 ;
     RECT  28.7 406.04 31.58 409.6 ;
     RECT  30.62 465.26 31.78 468.4 ;
     RECT  31.58 406.04 33.02 410.02 ;
     RECT  33.02 402.68 33.5 410.02 ;
     RECT  28.7 527 33.5 531.4 ;
     RECT  33.5 526.16 33.7 531.4 ;
     RECT  33.5 396.38 33.98 410.02 ;
     RECT  33.5 292.22 34.18 292.42 ;
     RECT  34.46 353.96 34.94 354.16 ;
     RECT  31.58 488.78 35.14 488.98 ;
     RECT  34.94 352.7 36.1 354.16 ;
     RECT  33.98 396.38 36.1 417.58 ;
     RECT  34.94 552.62 36.38 552.82 ;
     RECT  36.1 353.12 36.58 354.16 ;
     RECT  33.98 387.56 37.06 387.76 ;
     RECT  36.1 396.38 37.34 410.02 ;
     RECT  33.7 526.16 37.34 530.56 ;
     RECT  36.58 353.12 37.54 353.32 ;
     RECT  33.5 464.84 37.54 465.04 ;
     RECT  38.3 374.96 39.74 375.16 ;
     RECT  31.1 479.12 40.22 479.32 ;
     RECT  37.34 391.34 42.34 410.02 ;
     RECT  36.38 550.1 42.34 552.82 ;
     RECT  40.22 479.12 42.82 480.58 ;
     RECT  37.34 524.9 42.82 530.56 ;
     RECT  39.74 281.72 43.1 281.92 ;
     RECT  42.62 455.6 43.1 455.8 ;
     RECT  36.86 266.18 43.58 266.38 ;
     RECT  43.1 279.2 43.58 281.92 ;
     RECT  43.1 477.86 44.06 478.06 ;
     RECT  40.22 568.58 44.06 568.78 ;
     RECT  44.06 468.2 44.54 468.4 ;
     RECT  44.06 477.02 44.54 478.06 ;
     RECT  36.38 440.9 45.02 441.1 ;
     RECT  43.1 451.4 45.02 455.8 ;
     RECT  43.58 263.24 45.22 266.38 ;
     RECT  42.62 300.62 45.22 300.82 ;
     RECT  39.74 374.96 45.5 382.3 ;
     RECT  42.34 391.34 45.5 406.24 ;
     RECT  42.14 500.54 45.5 500.74 ;
     RECT  42.82 530.36 45.5 530.56 ;
     RECT  45.02 440.9 45.7 455.8 ;
     RECT  45.5 530.36 46.18 538.54 ;
     RECT  45.22 264.08 46.66 266.38 ;
     RECT  45.5 374.96 46.66 406.24 ;
     RECT  44.54 468.2 47.14 478.06 ;
     RECT  45.5 500.54 47.42 504.52 ;
     RECT  46.94 539.6 48.1 539.8 ;
     RECT  44.06 568.58 48.1 569.62 ;
     RECT  43.58 279.2 49.54 284.86 ;
     RECT  47.14 471.14 49.54 478.06 ;
     RECT  47.42 496.76 49.54 504.52 ;
     RECT  48.38 424.94 50.02 425.14 ;
     RECT  47.9 338 50.3 338.2 ;
     RECT  46.18 530.36 50.5 530.56 ;
     RECT  42.34 552.62 50.5 552.82 ;
     RECT  48.1 568.58 50.5 568.78 ;
     RECT  46.94 586.22 50.5 586.42 ;
     RECT  50.3 368.66 50.78 368.86 ;
     RECT  49.54 496.76 50.78 497.38 ;
     RECT  50.3 509.78 50.78 509.98 ;
     RECT  47.9 519.02 50.78 519.22 ;
     RECT  50.78 489.2 51.26 497.38 ;
     RECT  50.3 337.16 51.46 338.2 ;
     RECT  45.7 448.04 51.46 455.8 ;
     RECT  51.26 478.28 51.46 497.38 ;
     RECT  50.78 509.78 51.46 519.22 ;
     RECT  46.66 266.18 51.74 266.38 ;
     RECT  50.78 363.62 51.74 368.86 ;
     RECT  51.46 455.6 51.74 455.8 ;
     RECT  51.46 511.88 51.74 519.22 ;
     RECT  51.74 266.18 51.94 270.16 ;
     RECT  51.74 455.6 51.94 456.64 ;
     RECT  51.46 496.76 51.94 497.38 ;
     RECT  46.66 380.84 52.22 406.24 ;
     RECT  49.54 279.2 52.42 281.08 ;
     RECT  52.22 380.84 52.42 409.18 ;
     RECT  52.42 380.84 52.9 389.44 ;
     RECT  51.94 269.96 53.38 270.16 ;
     RECT  51.94 497.18 53.38 497.38 ;
     RECT  50.3 298.94 54.34 300.4 ;
     RECT  51.74 357.74 54.62 368.86 ;
     RECT  54.34 300.2 55.1 300.4 ;
     RECT  54.62 357.32 55.1 368.86 ;
     RECT  53.18 341.78 55.3 341.98 ;
     RECT  33.98 323.3 55.58 323.5 ;
     RECT  55.1 357.32 55.58 372.22 ;
     RECT  52.9 380.84 55.58 386.92 ;
     RECT  50.3 425.78 55.58 425.98 ;
     RECT  54.62 602.6 55.58 602.8 ;
     RECT  55.1 300.2 55.78 307.54 ;
     RECT  51.46 478.28 55.78 485.2 ;
     RECT  52.42 279.2 56.06 280.24 ;
     RECT  55.78 478.28 56.26 478.48 ;
     RECT  52.7 251.48 57.02 251.68 ;
     RECT  55.58 598.4 57.22 602.8 ;
     RECT  57.02 244.34 57.7 251.68 ;
     RECT  56.06 278.36 57.7 280.24 ;
     RECT  57.98 470.72 58.46 470.92 ;
     RECT  56.54 557.24 58.66 557.44 ;
     RECT  55.58 319.52 58.94 323.5 ;
     RECT  52.42 398.48 58.94 409.18 ;
     RECT  58.94 398.48 59.62 410.02 ;
     RECT  55.58 357.32 60.1 386.92 ;
     RECT  57.22 598.4 60.58 599.86 ;
     RECT  55.78 307.34 61.34 307.54 ;
     RECT  58.94 318.26 61.34 323.5 ;
     RECT  51.94 456.44 61.34 456.64 ;
     RECT  60.1 357.74 61.54 386.92 ;
     RECT  61.34 448.04 62.3 456.64 ;
     RECT  58.46 466.52 62.3 470.92 ;
     RECT  60.58 598.4 62.5 599.44 ;
     RECT  57.7 278.36 62.98 279.4 ;
     RECT  61.54 357.74 62.98 372.22 ;
     RECT  51.74 511.88 62.98 527.62 ;
     RECT  57.98 547.16 62.98 547.36 ;
     RECT  62.3 344.72 63.46 344.92 ;
     RECT  55.58 425.78 63.74 428.08 ;
     RECT  63.26 505.16 63.74 505.36 ;
     RECT  59.62 409.82 63.94 410.02 ;
     RECT  61.54 382.94 64.42 386.92 ;
     RECT  62.3 448.04 66.14 470.92 ;
     RECT  64.42 386.72 66.62 386.92 ;
     RECT  59.62 398.48 66.62 400.36 ;
     RECT  61.34 307.34 67.1 323.5 ;
     RECT  62.98 517.76 67.78 527.62 ;
     RECT  66.14 259.04 68.06 259.24 ;
     RECT  67.1 591.68 68.26 591.88 ;
     RECT  63.74 420.74 68.54 428.08 ;
     RECT  67.1 300.62 68.74 323.5 ;
     RECT  67.78 517.76 68.74 525.52 ;
     RECT  64.7 546.74 69.02 546.94 ;
     RECT  68.54 413.6 69.22 436.48 ;
     RECT  68.74 518.18 69.22 525.52 ;
     RECT  69.02 541.28 69.22 546.94 ;
     RECT  68.74 300.62 69.98 307.54 ;
     RECT  69.22 413.6 70.18 428.5 ;
     RECT  69.22 518.6 70.18 525.52 ;
     RECT  66.14 448.04 70.46 472.6 ;
     RECT  62.98 359.42 70.94 372.22 ;
     RECT  68.54 572.78 71.9 572.98 ;
     RECT  70.46 440.48 72.38 472.6 ;
     RECT  66.62 386.72 72.86 400.36 ;
     RECT  72.38 440.48 73.34 474.28 ;
     RECT  57.7 244.34 73.82 244.54 ;
     RECT  70.94 359.42 73.82 372.64 ;
     RECT  71.9 572.78 74.02 576.76 ;
     RECT  63.74 504.74 74.3 505.36 ;
     RECT  72.86 383.36 75.26 402.46 ;
     RECT  69.98 299.36 75.46 307.54 ;
     RECT  70.18 420.74 75.46 428.5 ;
     RECT  74.3 496.34 75.46 505.36 ;
     RECT  74.3 339.68 75.94 339.88 ;
     RECT  73.82 239.72 76.9 244.54 ;
     RECT  76.9 244.34 77.38 244.54 ;
     RECT  70.18 521.12 77.38 525.52 ;
     RECT  73.34 440.48 77.86 478.48 ;
     RECT  77.38 523.22 77.86 525.52 ;
     RECT  75.26 383.36 79.1 410.86 ;
     RECT  75.46 420.74 79.1 428.08 ;
     RECT  77.86 447.2 79.1 478.48 ;
     RECT  77.86 523.22 79.3 523.42 ;
     RECT  79.1 289.28 79.58 289.48 ;
     RECT  75.46 299.36 79.58 302.08 ;
     RECT  68.74 319.94 79.58 323.5 ;
     RECT  79.1 447.2 79.78 481.84 ;
     RECT  62.98 279.2 81.5 279.4 ;
     RECT  79.58 289.28 81.5 302.08 ;
     RECT  73.82 358.16 81.5 372.64 ;
     RECT  81.5 357.32 81.7 372.64 ;
     RECT  81.7 357.32 81.98 371.38 ;
     RECT  79.78 466.1 82.46 481.84 ;
     RECT  69.22 541.28 82.46 541.48 ;
     RECT  79.58 314.48 82.94 328.54 ;
     RECT  77.66 345.56 83.14 345.76 ;
     RECT  81.5 279.2 83.62 302.08 ;
     RECT  82.94 314.48 83.62 334.84 ;
     RECT  82.46 466.1 83.62 486.88 ;
     RECT  83.62 316.16 84.58 334.84 ;
     RECT  79.1 383.36 85.34 428.08 ;
     RECT  83.62 289.28 85.54 302.08 ;
     RECT  82.46 541.28 85.82 541.9 ;
     RECT  68.06 259.04 86.5 266.8 ;
     RECT  83.62 466.1 86.5 470.92 ;
     RECT  75.46 504.74 86.78 505.36 ;
     RECT  83.62 481.64 86.98 486.88 ;
     RECT  81.98 356.48 88.22 371.38 ;
     RECT  79.78 447.2 88.22 456.64 ;
     RECT  86.78 503.9 88.42 505.36 ;
     RECT  85.54 296.42 88.9 302.08 ;
     RECT  88.42 505.16 89.38 505.36 ;
     RECT  85.34 383.36 89.66 433.12 ;
     RECT  88.22 447.2 89.66 457.48 ;
     RECT  88.9 296.84 89.86 302.08 ;
     RECT  89.66 383.36 89.86 457.48 ;
     RECT  89.86 296.84 90.82 297.46 ;
     RECT  89.86 383.36 91.3 456.64 ;
     RECT  74.02 572.78 92.06 572.98 ;
     RECT  88.22 353.12 92.26 371.38 ;
     RECT  86.5 466.1 93.5 467.14 ;
     RECT  92.26 353.12 93.7 370.96 ;
     RECT  91.3 383.36 93.7 394.06 ;
     RECT  84.58 317.84 94.18 334.84 ;
     RECT  93.7 353.12 94.18 360.88 ;
     RECT  91.3 427.88 94.18 439 ;
     RECT  94.18 327.08 94.94 334.84 ;
     RECT  92.06 568.58 94.94 572.98 ;
     RECT  92.54 251.06 95.14 251.26 ;
     RECT  91.3 447.62 95.14 456.64 ;
     RECT  93.5 465.26 95.42 467.14 ;
     RECT  93.7 383.36 96.1 387.34 ;
     RECT  94.18 432.92 96.1 439 ;
     RECT  93.02 599.24 96.86 599.44 ;
     RECT  94.18 360.26 97.06 360.88 ;
     RECT  96.1 383.36 97.06 385.66 ;
     RECT  90.82 297.26 97.54 297.46 ;
     RECT  96.1 438.8 97.54 439 ;
     RECT  79.1 149.42 98.02 149.62 ;
     RECT  97.06 360.68 98.02 360.88 ;
     RECT  95.42 465.26 98.3 474.7 ;
     RECT  91.3 402.68 98.5 413.38 ;
     RECT  94.94 568.58 98.78 576.76 ;
     RECT  94.94 327.08 98.98 343.24 ;
     RECT  98.3 459.8 99.46 474.7 ;
     RECT  98.98 327.5 100.7 343.24 ;
     RECT  86.5 263.24 100.9 266.8 ;
     RECT  94.18 317.84 100.9 318.46 ;
     RECT  96.86 599.24 100.9 601.96 ;
     RECT  95.14 447.62 101.38 448.24 ;
     RECT  98.5 413.18 102.14 413.38 ;
     RECT  101.18 523.64 102.14 523.84 ;
     RECT  99.46 462.32 103.58 474.7 ;
     RECT  86.98 486.68 103.58 486.88 ;
     RECT  102.14 413.18 104.26 420.94 ;
     RECT  102.14 520.28 104.54 523.84 ;
     RECT  85.82 539.18 105.5 541.9 ;
     RECT  103.58 462.32 106.18 486.88 ;
     RECT  95.42 550.52 106.46 554.08 ;
     RECT  98.78 568.16 106.46 576.76 ;
     RECT  104.54 520.28 106.94 526.78 ;
     RECT  105.5 535.82 106.94 541.9 ;
     RECT  106.46 550.52 106.94 576.76 ;
     RECT  46.46 219.56 107.42 219.76 ;
     RECT  97.34 504.32 107.42 504.52 ;
     RECT  106.94 519.02 107.42 576.76 ;
     RECT  100.9 600.5 107.42 601.96 ;
     RECT  106.18 462.32 107.62 473.86 ;
     RECT  100.9 318.26 107.9 318.46 ;
     RECT  100.7 327.5 107.9 348.28 ;
     RECT  106.18 486.68 107.9 486.88 ;
     RECT  107.42 504.32 108.86 576.76 ;
     RECT  107.9 318.26 109.34 348.28 ;
     RECT  93.7 370.76 109.34 370.96 ;
     RECT  107.42 600.5 109.34 610.36 ;
     RECT  97.06 385.46 109.82 385.66 ;
     RECT  109.34 600.5 109.82 615.4 ;
     RECT  76.22 111.62 110.5 111.82 ;
     RECT  109.34 318.26 110.5 349.54 ;
     RECT  107.62 468.62 110.5 473.86 ;
     RECT  109.34 370.76 111.26 372.64 ;
     RECT  108.38 430.82 111.26 431.02 ;
     RECT  83.62 279.2 111.74 279.4 ;
     RECT  100.7 288.86 111.74 289.06 ;
     RECT  110.5 318.26 111.74 348.28 ;
     RECT  111.26 430.82 112.7 432.7 ;
     RECT  102.62 442.58 112.7 442.78 ;
     RECT  112.7 430.82 112.9 442.78 ;
     RECT  109.82 600.5 112.9 617.92 ;
     RECT  112.9 440.48 113.38 442.78 ;
     RECT  111.74 317 113.66 348.28 ;
     RECT  104.26 419.06 113.66 420.94 ;
     RECT  112.9 430.82 113.66 431.02 ;
     RECT  113.66 419.06 113.86 431.02 ;
     RECT  112.9 600.5 113.86 615.4 ;
     RECT  111.26 368.24 114.14 372.64 ;
     RECT  109.82 385.46 114.14 389.02 ;
     RECT  113.38 442.58 114.14 442.78 ;
     RECT  108.86 497.6 114.82 576.76 ;
     RECT  108.38 587.9 115.1 588.1 ;
     RECT  113.86 600.5 115.3 610.36 ;
     RECT  111.74 279.2 115.58 289.06 ;
     RECT  115.58 279.2 116.54 289.48 ;
     RECT  114.14 368.24 117.02 389.02 ;
     RECT  110.5 469.04 117.02 473.86 ;
     RECT  116.54 279.2 117.5 289.9 ;
     RECT  115.1 246.86 117.98 247.06 ;
     RECT  117.02 469.04 117.98 474.7 ;
     RECT  107.9 486.68 117.98 487.3 ;
     RECT  114.82 497.6 117.98 575.92 ;
     RECT  117.5 277.94 118.46 289.9 ;
     RECT  106.94 300.62 118.46 300.82 ;
     RECT  113.66 315.74 118.46 348.28 ;
     RECT  117.02 361.52 119.62 389.02 ;
     RECT  117.98 469.04 119.9 575.92 ;
     RECT  117.98 246.86 122.02 251.68 ;
     RECT  119.9 468.2 122.02 575.92 ;
     RECT  122.02 468.2 122.3 475.54 ;
     RECT  118.46 277.94 122.78 348.28 ;
     RECT  114.14 442.58 122.78 444.04 ;
     RECT  120.86 454.76 122.78 454.96 ;
     RECT  115.3 600.5 122.98 600.7 ;
     RECT  121.82 647.54 122.98 647.74 ;
     RECT  122.78 272.06 123.26 348.28 ;
     RECT  117.5 400.16 123.26 400.36 ;
     RECT  122.3 467.78 123.74 475.54 ;
     RECT  122.02 486.68 123.94 575.92 ;
     RECT  123.26 400.16 124.22 402.88 ;
     RECT  115.1 584.54 124.22 588.1 ;
     RECT  115.3 610.16 124.22 610.36 ;
     RECT  124.22 400.16 124.7 406.66 ;
     RECT  113.86 419.06 124.7 427.24 ;
     RECT  123.26 266.6 125.38 348.28 ;
     RECT  125.38 307.76 126.34 331.06 ;
     RECT  122.78 442.58 126.34 454.96 ;
     RECT  119.62 368.24 127.1 389.02 ;
     RECT  124.7 400.16 127.1 427.24 ;
     RECT  124.22 610.16 127.3 613.3 ;
     RECT  126.34 307.76 128.26 307.96 ;
     RECT  125.38 342.62 129.02 348.28 ;
     RECT  126.34 447.2 129.02 454.96 ;
     RECT  123.74 464.42 129.02 475.54 ;
     RECT  127.1 368.24 129.7 427.24 ;
     RECT  129.7 368.24 130.46 403.72 ;
     RECT  129.02 447.2 130.46 475.54 ;
     RECT  123.94 486.68 130.46 572.56 ;
     RECT  125.38 266.6 131.14 297.88 ;
     RECT  131.14 266.6 131.62 287.38 ;
     RECT  129.02 342.62 131.9 352.9 ;
     RECT  131.9 342.62 133.06 353.32 ;
     RECT  130.46 367.82 133.34 403.72 ;
     RECT  127.3 610.16 133.34 610.36 ;
     RECT  122.02 247.28 133.54 251.68 ;
     RECT  124.22 584.12 133.54 588.1 ;
     RECT  129.5 651.74 133.54 651.94 ;
     RECT  133.34 367.4 133.82 403.72 ;
     RECT  131.14 296.84 134.02 297.88 ;
     RECT  133.82 365.72 134.02 403.72 ;
     RECT  133.34 609.32 134.02 610.36 ;
     RECT  130.46 447.2 134.5 572.56 ;
     RECT  133.06 342.62 134.78 352.9 ;
     RECT  129.7 413.6 135.26 427.24 ;
     RECT  127.1 437.96 135.26 438.58 ;
     RECT  135.74 195.62 136.42 195.82 ;
     RECT  133.54 248.12 136.42 251.68 ;
     RECT  131.62 266.6 136.9 279.4 ;
     RECT  134.78 307.34 136.9 307.54 ;
     RECT  126.34 316.58 136.9 331.06 ;
     RECT  134.02 366.56 136.9 403.72 ;
     RECT  136.9 317 137.38 331.06 ;
     RECT  137.38 317 137.86 317.2 ;
     RECT  135.26 413.6 138.14 438.58 ;
     RECT  134.5 447.2 138.14 475.54 ;
     RECT  107.42 219.56 138.34 225.22 ;
     RECT  136.7 629.48 138.62 629.68 ;
     RECT  134.02 296.84 139.78 297.04 ;
     RECT  137.38 327.5 140.26 331.06 ;
     RECT  136.7 652.16 140.54 652.36 ;
     RECT  138.62 628.64 141.22 629.68 ;
     RECT  140.54 593.78 141.5 593.98 ;
     RECT  134.78 341.78 142.46 352.9 ;
     RECT  133.54 584.12 142.94 584.32 ;
     RECT  141.5 593.78 142.94 595.24 ;
     RECT  136.42 248.12 143.14 251.26 ;
     RECT  138.14 413.6 143.42 475.54 ;
     RECT  142.46 341.78 143.9 357.52 ;
     RECT  143.42 413.18 143.9 475.54 ;
     RECT  134.5 486.68 143.9 572.56 ;
     RECT  138.34 219.56 144.38 219.76 ;
     RECT  140.54 652.16 144.86 656.56 ;
     RECT  141.22 628.64 146.02 628.84 ;
     RECT  143.9 334.64 146.78 357.52 ;
     RECT  144.86 647.54 146.98 656.56 ;
     RECT  144.38 217.04 147.46 219.76 ;
     RECT  146.98 647.54 147.94 655.72 ;
     RECT  136.9 266.6 148.22 266.8 ;
     RECT  146.78 334.64 148.22 357.94 ;
     RECT  136.9 367.82 148.22 403.72 ;
     RECT  136.9 279.2 149.18 279.4 ;
     RECT  148.7 288.86 149.18 289.06 ;
     RECT  142.94 584.12 150.34 595.24 ;
     RECT  148.22 334.64 150.62 403.72 ;
     RECT  143.14 248.12 150.82 248.32 ;
     RECT  148.22 266.6 151.1 269.74 ;
     RECT  149.18 279.2 151.1 289.06 ;
     RECT  143.9 413.18 151.1 572.56 ;
     RECT  150.34 584.12 151.1 586.84 ;
     RECT  151.1 264.08 151.58 289.06 ;
     RECT  150.62 334.22 151.58 403.72 ;
     RECT  151.1 413.18 151.58 586.84 ;
     RECT  150.62 609.32 151.58 609.52 ;
     RECT  151.58 264.08 151.78 290.74 ;
     RECT  151.58 334.22 152.26 586.84 ;
     RECT  152.06 167.48 152.74 167.68 ;
     RECT  151.58 597.98 152.74 609.52 ;
     RECT  152.06 243.92 153.02 247.48 ;
     RECT  150.62 305.24 153.02 305.44 ;
     RECT  151.1 196.88 153.5 197.08 ;
     RECT  153.02 323.3 153.5 323.5 ;
     RECT  152.26 334.22 153.5 572.56 ;
     RECT  152.74 597.98 153.7 600.28 ;
     RECT  151.78 266.6 154.18 290.74 ;
     RECT  153.5 196.88 154.46 198.76 ;
     RECT  153.02 305.24 154.46 305.86 ;
     RECT  154.18 266.6 155.14 289.06 ;
     RECT  154.46 189.74 155.42 198.76 ;
     RECT  153.5 323.3 156.58 572.56 ;
     RECT  155.42 189.74 156.86 202.54 ;
     RECT  147.46 217.46 156.86 219.76 ;
     RECT  155.9 668.12 158.02 668.32 ;
     RECT  156.86 215.78 158.78 219.76 ;
     RECT  158.3 636.2 159.26 636.4 ;
     RECT  147.94 648.8 159.94 649 ;
     RECT  155.14 266.6 161.38 270.16 ;
     RECT  153.02 237.62 161.66 247.48 ;
     RECT  152.06 621.92 162.14 622.12 ;
     RECT  158.78 215.78 163.3 221.86 ;
     RECT  162.14 621.92 163.58 625.06 ;
     RECT  159.26 635.78 163.58 636.4 ;
     RECT  155.14 279.62 164.06 289.06 ;
     RECT  153.7 600.08 164.54 600.28 ;
     RECT  152.74 609.32 164.54 609.52 ;
     RECT  164.54 600.08 165.02 609.52 ;
     RECT  165.02 600.08 165.5 610.36 ;
     RECT  163.58 621.92 165.5 636.4 ;
     RECT  161.38 268.28 165.98 270.16 ;
     RECT  164.06 279.2 165.98 289.06 ;
     RECT  156.58 323.3 165.98 452.02 ;
     RECT  156.86 189.74 166.46 207.16 ;
     RECT  163.3 215.78 166.46 219.76 ;
     RECT  166.46 189.74 166.94 219.76 ;
     RECT  165.5 600.08 167.14 636.4 ;
     RECT  165.98 268.28 167.9 289.06 ;
     RECT  156.58 464.42 168.38 572.56 ;
     RECT  165.98 322.46 168.86 452.02 ;
     RECT  168.38 461.9 168.86 572.56 ;
     RECT  162.14 647.96 169.06 648.16 ;
     RECT  167.9 268.28 169.34 289.9 ;
     RECT  154.46 303.14 169.34 305.86 ;
     RECT  154.46 694.58 169.34 694.78 ;
     RECT  165.5 103.64 169.54 103.84 ;
     RECT  163.1 259.04 169.54 259.24 ;
     RECT  168.38 133.46 169.82 133.66 ;
     RECT  168.86 322.46 170.3 572.56 ;
     RECT  152.26 584.12 170.3 586.84 ;
     RECT  161.66 232.16 170.5 247.48 ;
     RECT  170.3 322.46 170.5 586.84 ;
     RECT  170.5 232.16 170.78 244.96 ;
     RECT  169.34 268.28 170.78 305.86 ;
     RECT  170.5 322.46 171.26 475.54 ;
     RECT  171.26 318.26 171.46 475.54 ;
     RECT  166.94 189.32 172.22 219.76 ;
     RECT  170.78 228.8 172.22 244.96 ;
     RECT  172.22 189.32 172.42 244.96 ;
     RECT  169.82 133.46 172.9 140.38 ;
     RECT  172.42 189.32 173.66 202.96 ;
     RECT  172.42 214.1 173.86 244.96 ;
     RECT  173.86 214.1 174.82 229 ;
     RECT  173.86 243.5 176.26 244.96 ;
     RECT  170.78 262.82 177.5 305.86 ;
     RECT  171.46 318.26 177.5 370.12 ;
     RECT  177.5 262.82 177.7 370.12 ;
     RECT  172.9 137.66 177.98 140.38 ;
     RECT  177.7 262.82 177.98 338.2 ;
     RECT  167.14 621.92 178.46 636.4 ;
     RECT  171.46 378.74 178.94 475.54 ;
     RECT  170.5 485.84 178.94 586.84 ;
     RECT  165.02 172.52 179.42 172.72 ;
     RECT  167.14 600.08 179.42 610.36 ;
     RECT  178.46 621.5 179.42 636.4 ;
     RECT  177.7 349.76 179.9 370.12 ;
     RECT  178.94 378.74 179.9 586.84 ;
     RECT  179.42 600.08 180.38 636.4 ;
     RECT  180.38 600.08 181.82 640.18 ;
     RECT  179.9 349.76 182.02 586.84 ;
     RECT  177.98 137.66 182.5 142.06 ;
     RECT  173.66 186.38 182.98 202.96 ;
     RECT  174.82 214.1 183.26 219.76 ;
     RECT  179.42 168.32 183.46 172.72 ;
     RECT  177.98 259.88 183.94 338.2 ;
     RECT  181.82 600.08 184.22 645.22 ;
     RECT  182.98 186.8 184.42 202.96 ;
     RECT  185.66 156.14 186.62 156.34 ;
     RECT  183.46 168.32 186.62 171.46 ;
     RECT  182.5 137.66 186.82 140.38 ;
     RECT  184.22 599.24 186.82 645.22 ;
     RECT  186.62 151.52 188.06 156.34 ;
     RECT  186.62 164.96 188.06 171.46 ;
     RECT  188.06 151.52 188.26 171.46 ;
     RECT  176.26 244.76 188.74 244.96 ;
     RECT  182.02 351.02 188.74 586.84 ;
     RECT  186.82 600.08 189.22 645.22 ;
     RECT  169.34 694.58 190.46 697.72 ;
     RECT  189.22 600.08 190.66 644.38 ;
     RECT  190.46 689.12 191.42 697.72 ;
     RECT  183.26 213.68 191.9 219.76 ;
     RECT  190.66 610.16 192.1 639.76 ;
     RECT  192.1 610.16 192.58 628.42 ;
     RECT  183.94 269.54 193.06 338.2 ;
     RECT  190.66 600.08 193.54 600.28 ;
     RECT  184.42 186.8 193.82 200.86 ;
     RECT  191.9 213.26 193.82 219.76 ;
     RECT  183.94 259.88 193.82 260.08 ;
     RECT  188.26 164.12 194.3 171.46 ;
     RECT  193.82 186.8 194.3 219.76 ;
     RECT  192.58 610.16 194.5 610.36 ;
     RECT  186.82 140.18 195.74 140.38 ;
     RECT  188.26 151.52 195.74 151.72 ;
     RECT  194.3 164.12 195.74 219.76 ;
     RECT  174.82 228.8 195.74 229 ;
     RECT  195.74 140.18 196.7 151.72 ;
     RECT  195.74 164.12 196.9 229 ;
     RECT  196.9 164.12 197.38 200.86 ;
     RECT  193.06 269.54 197.38 315.1 ;
     RECT  188.74 380 197.38 586.84 ;
     RECT  197.38 164.12 197.86 169.78 ;
     RECT  197.38 314.9 199.3 315.1 ;
     RECT  188.74 351.02 199.3 370.12 ;
     RECT  196.7 140.18 199.58 152.98 ;
     RECT  197.86 164.12 199.58 168.94 ;
     RECT  197.38 380 200.74 575.08 ;
     RECT  192.1 639.56 200.74 639.76 ;
     RECT  193.82 251.48 201.02 260.08 ;
     RECT  196.9 212.42 201.5 229 ;
     RECT  193.06 324.98 201.5 338.2 ;
     RECT  199.3 351.02 201.5 353.32 ;
     RECT  192.58 621.92 201.5 628.42 ;
     RECT  201.5 324.98 201.98 353.32 ;
     RECT  201.5 621.92 201.98 629.26 ;
     RECT  197.66 652.16 202.66 652.36 ;
     RECT  199.3 363.62 202.94 370.12 ;
     RECT  200.74 380 202.94 572.14 ;
     RECT  199.58 140.18 203.9 168.94 ;
     RECT  203.9 610.16 204.38 610.36 ;
     RECT  201.5 212.42 204.86 232.36 ;
     RECT  204.38 602.6 204.86 610.36 ;
     RECT  204.86 212.42 205.34 239.92 ;
     RECT  201.02 249.38 205.34 260.08 ;
     RECT  197.38 269.54 205.34 305.86 ;
     RECT  204.86 602.18 205.82 610.78 ;
     RECT  201.98 621.92 205.82 629.68 ;
     RECT  197.38 584.12 207.26 586.84 ;
     RECT  197.38 178.4 207.46 200.86 ;
     RECT  203.9 138.08 207.74 168.94 ;
     RECT  207.46 197.3 207.74 200.86 ;
     RECT  205.34 212.42 207.74 305.86 ;
     RECT  201.98 315.32 208.22 353.32 ;
     RECT  207.74 197.3 208.7 305.86 ;
     RECT  208.22 314.9 208.7 353.32 ;
     RECT  202.94 363.62 208.7 572.14 ;
     RECT  208.7 197.3 209.18 572.14 ;
     RECT  207.26 584.12 209.18 589.78 ;
     RECT  205.82 602.18 209.18 629.68 ;
     RECT  209.18 197.3 209.66 572.56 ;
     RECT  209.18 584.12 209.66 629.68 ;
     RECT  207.46 178.4 210.34 187.84 ;
     RECT  209.18 652.58 210.62 652.78 ;
     RECT  209.66 197.3 211.1 629.68 ;
     RECT  210.62 652.58 213.02 657.4 ;
     RECT  213.02 652.58 213.98 664.12 ;
     RECT  211.1 197.3 215.14 635.98 ;
     RECT  207.74 130.52 216.86 168.94 ;
     RECT  210.34 178.4 216.86 187.42 ;
     RECT  215.14 353.12 216.86 635.98 ;
     RECT  215.14 197.3 217.34 341.56 ;
     RECT  216.86 353.12 217.82 638.08 ;
     RECT  216.86 130.52 218.5 187.42 ;
     RECT  217.34 196.46 218.5 341.56 ;
     RECT  218.5 196.46 219.94 234.88 ;
     RECT  218.5 243.5 220.42 341.56 ;
     RECT  217.82 353.12 220.7 640.18 ;
     RECT  220.7 353.12 221.18 640.6 ;
     RECT  213.98 652.16 221.18 664.12 ;
     RECT  218.5 130.52 222.82 187 ;
     RECT  221.18 353.12 222.82 664.12 ;
     RECT  219.94 196.46 223.78 232.36 ;
     RECT  222.82 582.86 223.78 664.12 ;
     RECT  222.82 130.52 224.74 186.58 ;
     RECT  223.78 198.14 226.18 232.36 ;
     RECT  224.74 130.52 226.66 161.38 ;
     RECT  222.82 353.12 226.66 572.56 ;
     RECT  224.74 171.26 228.58 186.58 ;
     RECT  226.18 198.14 229.06 224.38 ;
     RECT  226.66 353.12 229.54 560.38 ;
     RECT  229.06 201.08 230.5 224.38 ;
     RECT  220.42 243.5 230.78 255.04 ;
     RECT  220.42 267.02 230.78 341.56 ;
     RECT  230.78 243.5 230.98 341.56 ;
     RECT  229.54 363.62 230.98 560.38 ;
     RECT  223.78 582.86 231.26 600.28 ;
     RECT  230.98 243.5 231.94 258.82 ;
     RECT  231.26 582.44 232.22 600.28 ;
     RECT  223.78 609.74 232.22 664.12 ;
     RECT  228.58 171.26 232.42 179.86 ;
     RECT  230.5 205.7 232.42 224.38 ;
     RECT  231.94 248.96 232.9 258.82 ;
     RECT  230.98 363.62 232.9 550.72 ;
     RECT  226.66 130.52 233.38 160.96 ;
     RECT  232.42 171.26 233.86 179.44 ;
     RECT  230.98 559.76 236.06 560.38 ;
     RECT  226.66 572.36 236.06 572.56 ;
     RECT  232.42 213.68 236.26 224.38 ;
     RECT  233.38 156.56 237.5 160.96 ;
     RECT  233.86 171.26 237.5 175.24 ;
     RECT  230.98 269.54 237.7 341.56 ;
     RECT  236.06 559.76 237.7 572.56 ;
     RECT  237.7 314.9 238.18 341.56 ;
     RECT  237.7 572.36 239.42 572.56 ;
     RECT  232.22 582.44 239.42 664.12 ;
     RECT  237.5 156.56 240.58 175.24 ;
     RECT  229.54 353.12 240.86 353.74 ;
     RECT  232.9 363.62 240.86 371.8 ;
     RECT  232.9 383.78 241.34 550.72 ;
     RECT  237.7 559.76 241.34 560.38 ;
     RECT  240.86 353.12 241.54 371.8 ;
     RECT  239.42 572.36 241.54 664.12 ;
     RECT  161.66 673.16 241.82 673.36 ;
     RECT  191.42 689.12 241.82 698.98 ;
     RECT  237.7 269.54 242.02 305.86 ;
     RECT  241.54 363.62 242.3 371.8 ;
     RECT  241.54 584.12 242.3 664.12 ;
     RECT  241.82 673.16 242.3 698.98 ;
     RECT  240.58 160.76 243.46 175.24 ;
     RECT  242.3 584.12 243.46 698.98 ;
     RECT  243.46 163.7 244.7 175.24 ;
     RECT  242.02 285.08 244.9 305.86 ;
     RECT  243.46 584.12 244.9 663.28 ;
     RECT  241.54 353.12 245.38 354.16 ;
     RECT  241.34 383.78 245.38 560.38 ;
     RECT  244.7 163.7 246.14 183.64 ;
     RECT  232.9 251.9 246.14 258.82 ;
     RECT  242.02 269.54 246.14 270.16 ;
     RECT  236.26 224.18 246.82 224.38 ;
     RECT  238.18 316.16 247.1 341.56 ;
     RECT  244.9 288.86 247.3 305.86 ;
     RECT  244.9 584.12 247.3 630.52 ;
     RECT  244.9 639.56 247.3 663.28 ;
     RECT  247.1 316.16 247.78 342.82 ;
     RECT  246.14 251.9 248.26 270.16 ;
     RECT  247.3 642.08 248.74 663.28 ;
     RECT  247.3 288.86 249.22 292.42 ;
     RECT  247.78 318.68 249.7 342.82 ;
     RECT  246.14 163.7 250.66 191.62 ;
     RECT  247.58 228.8 250.66 229 ;
     RECT  249.22 291.38 250.66 292.42 ;
     RECT  245.38 385.04 250.66 560.38 ;
     RECT  248.26 259.46 251.14 270.16 ;
     RECT  247.3 617.72 251.14 630.52 ;
     RECT  245.38 353.54 251.62 354.16 ;
     RECT  242.3 363.62 251.62 372.22 ;
     RECT  250.66 163.7 252.1 175.24 ;
     RECT  250.66 191.42 252.1 191.62 ;
     RECT  249.7 320.36 252.1 342.82 ;
     RECT  252.1 168.32 253.06 168.52 ;
     RECT  251.62 363.62 253.34 368.86 ;
     RECT  252.1 320.36 253.54 334.84 ;
     RECT  241.54 572.36 254.3 572.56 ;
     RECT  247.3 584.12 254.3 608.68 ;
     RECT  254.3 572.36 254.78 608.68 ;
     RECT  253.34 355.22 254.98 368.86 ;
     RECT  233.38 130.52 255.46 147.52 ;
     RECT  255.46 138.08 255.94 147.52 ;
     RECT  255.94 138.08 256.42 138.28 ;
     RECT  250.66 385.04 256.7 550.72 ;
     RECT  251.14 617.72 256.7 629.68 ;
     RECT  248.74 642.08 256.7 660.76 ;
     RECT  251.14 259.46 256.9 259.66 ;
     RECT  254.78 561.86 257.66 608.68 ;
     RECT  256.7 617.3 257.66 629.68 ;
     RECT  256.7 638.72 257.86 660.76 ;
     RECT  256.7 382.1 260.06 550.72 ;
     RECT  257.66 561.86 260.06 629.68 ;
     RECT  251.14 269.54 260.26 270.16 ;
     RECT  260.06 382.1 261.98 629.68 ;
     RECT  257.86 638.72 261.98 660.34 ;
     RECT  261.98 382.1 262.66 660.34 ;
     RECT  253.54 321.2 263.9 334.84 ;
     RECT  262.66 382.1 263.9 659.92 ;
     RECT  260.26 269.54 265.06 269.74 ;
     RECT  263.9 321.2 265.06 342.4 ;
     RECT  247.3 304.4 266.02 305.86 ;
     RECT  265.06 321.2 269.86 334.84 ;
     RECT  255.94 147.32 270.34 147.52 ;
     RECT  269.86 334.64 270.82 334.84 ;
     RECT  266.02 304.4 271.3 304.6 ;
     RECT  269.86 321.2 271.78 321.4 ;
     RECT  250.66 292.22 272.54 292.42 ;
     RECT  254.98 359 272.54 368.86 ;
     RECT  263.9 381.68 272.54 659.92 ;
     RECT  272.54 381.22 273.02 659.92 ;
     RECT  272.54 292.22 276.1 298.26 ;
     RECT  275.9 339.64 276.38 339.84 ;
     RECT  277.82 173.74 278.3 173.94 ;
     RECT  276.38 339.64 279.74 342.36 ;
     RECT  279.74 313.6 280.22 313.8 ;
     RECT  279.26 226.24 280.7 226.44 ;
     RECT  276.86 142.66 282.62 142.86 ;
     RECT  270.62 154 282.62 154.2 ;
     RECT  281.66 272.44 282.62 272.64 ;
     RECT  279.74 334.18 282.62 342.36 ;
     RECT  280.7 226.24 283.78 228.96 ;
     RECT  280.22 311.5 284.06 313.8 ;
     RECT  282.14 282.52 284.54 282.72 ;
     RECT  282.62 142.66 284.74 154.2 ;
     RECT  282.62 327.88 284.74 342.36 ;
     RECT  282.62 269.08 285.02 272.64 ;
     RECT  273.02 381.22 285.5 663.7 ;
     RECT  284.54 282.52 285.98 286.92 ;
     RECT  276.1 298.06 285.98 298.26 ;
     RECT  270.62 203.56 286.18 203.76 ;
     RECT  285.98 282.52 286.46 298.26 ;
     RECT  284.06 309.4 286.46 313.8 ;
     RECT  286.46 282.52 287.42 315.06 ;
     RECT  284.74 335.44 287.42 342.36 ;
     RECT  272.54 354.34 287.42 368.86 ;
     RECT  285.5 380.38 287.42 663.7 ;
     RECT  281.66 131.74 288.1 131.94 ;
     RECT  284.74 142.66 288.38 143.28 ;
     RECT  285.02 267.4 288.38 272.64 ;
     RECT  288.38 266.98 289.34 272.64 ;
     RECT  284.74 154 289.54 154.2 ;
     RECT  289.34 266.56 289.54 272.64 ;
     RECT  287.42 282.52 289.54 318 ;
     RECT  287.9 222.46 290.02 222.66 ;
     RECT  287.42 335.44 290.02 663.7 ;
     RECT  287.9 211.96 290.3 212.16 ;
     RECT  289.54 286.72 290.5 318 ;
     RECT  290.5 303.94 290.78 318 ;
     RECT  290.5 286.72 290.98 294.48 ;
     RECT  290.98 294.28 292.42 294.48 ;
     RECT  290.78 303.94 293.18 320.52 ;
     RECT  290.02 335.44 293.18 659.5 ;
     RECT  293.18 303.94 293.38 659.5 ;
     RECT  290.78 160.72 294.82 162.18 ;
     RECT  278.3 173.74 294.82 174.78 ;
     RECT  290.3 211.96 297.22 218.46 ;
     RECT  289.54 266.98 297.98 272.64 ;
     RECT  288.38 135.52 299.14 143.28 ;
     RECT  293.38 303.94 299.42 368.86 ;
     RECT  297.98 266.98 300.58 275.58 ;
     RECT  299.42 286.3 300.58 286.5 ;
     RECT  300.58 266.98 300.86 269.28 ;
     RECT  293.38 377.44 300.86 659.5 ;
     RECT  243.46 673.16 300.86 698.98 ;
     RECT  288.38 109.06 301.06 109.26 ;
     RECT  299.42 203.56 301.82 203.76 ;
     RECT  300.86 266.56 302.5 269.28 ;
     RECT  275.9 244.72 303.46 244.92 ;
     RECT  294.82 161.14 304.22 162.18 ;
     RECT  301.34 131.74 304.42 131.94 ;
     RECT  296.06 232.54 305.38 232.74 ;
     RECT  301.82 197.68 305.86 203.76 ;
     RECT  299.42 297.64 306.34 368.86 ;
     RECT  304.22 154 306.62 162.18 ;
     RECT  306.34 334.6 306.82 368.86 ;
     RECT  297.98 177.1 308.74 177.3 ;
     RECT  306.34 297.64 309.22 320.52 ;
     RECT  306.82 335.86 309.22 368.86 ;
     RECT  300.86 377.44 309.7 698.98 ;
     RECT  305.86 197.68 310.94 202.92 ;
     RECT  297.22 218.26 311.14 218.46 ;
     RECT  309.22 337.12 311.14 368.86 ;
     RECT  309.7 377.44 311.14 377.64 ;
     RECT  306.62 154 312.1 165.12 ;
     RECT  309.22 298.06 312.58 320.52 ;
     RECT  312.58 303.94 313.54 320.52 ;
     RECT  311.14 359 313.54 368.86 ;
     RECT  313.54 359 314.02 366.34 ;
     RECT  312.1 156.52 314.5 165.12 ;
     RECT  314.02 363.62 314.98 366.34 ;
     RECT  313.54 304.36 315.94 320.52 ;
     RECT  309.7 386.3 315.94 698.98 ;
     RECT  314.98 364.04 316.42 366.34 ;
     RECT  310.94 195.58 316.9 202.92 ;
     RECT  315.94 306.46 316.9 320.52 ;
     RECT  314.5 164.92 317.66 165.12 ;
     RECT  316.9 195.58 317.86 195.78 ;
     RECT  316.9 308.98 317.86 320.52 ;
     RECT  311.14 337.12 317.86 348.66 ;
     RECT  302.5 269.08 318.62 269.28 ;
     RECT  318.62 260.68 321.5 269.28 ;
     RECT  320.06 237.16 321.98 237.36 ;
     RECT  317.66 287.56 321.98 287.76 ;
     RECT  321.5 260.26 322.46 269.28 ;
     RECT  321.5 377.44 322.46 377.64 ;
     RECT  317.66 164.92 322.94 168.9 ;
     RECT  321.98 233.8 323.42 237.36 ;
     RECT  322.94 157.78 323.62 176.88 ;
     RECT  322.46 377.44 325.54 381.42 ;
     RECT  320.06 214.48 326.78 214.68 ;
     RECT  322.46 259.84 326.78 274.74 ;
     RECT  321.98 287.56 326.78 291.54 ;
     RECT  326.78 259.84 326.98 291.54 ;
     RECT  316.42 366.14 327.46 366.34 ;
     RECT  318.62 101.5 328.42 101.7 ;
     RECT  326.98 260.26 328.9 291.54 ;
     RECT  323.42 226.24 329.18 237.36 ;
     RECT  317.86 308.98 329.18 312.96 ;
     RECT  329.18 308.98 329.38 313.38 ;
     RECT  329.18 226.24 330.14 241.14 ;
     RECT  326.78 214.06 330.62 214.68 ;
     RECT  330.14 226.24 330.62 241.56 ;
     RECT  330.62 214.06 332.06 241.56 ;
     RECT  328.9 260.68 332.26 291.54 ;
     RECT  323.62 172.9 332.54 176.88 ;
     RECT  322.46 135.1 333.7 135.3 ;
     RECT  323.62 157.78 333.98 161.76 ;
     RECT  333.98 151.06 334.46 161.76 ;
     RECT  317.86 339.64 334.46 348.66 ;
     RECT  332.06 214.06 335.62 247.44 ;
     RECT  334.46 150.22 335.9 161.76 ;
     RECT  332.54 172.9 336.58 184.86 ;
     RECT  329.38 308.98 337.34 309.6 ;
     RECT  332.06 369.88 337.34 370.08 ;
     RECT  325.54 381.22 337.34 381.42 ;
     RECT  332.26 264.04 338.5 291.54 ;
     RECT  337.34 362.74 338.98 370.08 ;
     RECT  337.34 305.2 339.26 309.6 ;
     RECT  333.98 324.1 339.26 324.3 ;
     RECT  337.34 381.22 339.46 381.84 ;
     RECT  336.58 176.68 339.94 184.86 ;
     RECT  339.94 176.68 341.38 176.88 ;
     RECT  334.46 335.44 343.1 348.66 ;
     RECT  335.9 138.88 343.3 161.76 ;
     RECT  338.5 264.04 343.78 288.18 ;
     RECT  335.62 214.06 344.54 234 ;
     RECT  338.98 369.88 344.74 370.08 ;
     RECT  343.3 143.08 346.46 161.76 ;
     RECT  346.46 143.08 346.66 165.96 ;
     RECT  344.54 205.24 346.94 205.44 ;
     RECT  344.54 214.06 346.94 236.94 ;
     RECT  315.94 392.6 346.94 698.98 ;
     RECT  339.74 195.58 347.14 195.78 ;
     RECT  343.78 283.36 347.9 288.18 ;
     RECT  343.78 264.04 348.38 271.38 ;
     RECT  348.38 262.78 348.86 271.38 ;
     RECT  339.26 305.2 349.06 324.3 ;
     RECT  339.46 381.22 349.34 381.42 ;
     RECT  346.94 392.56 349.34 698.98 ;
     RECT  348.86 262.36 349.82 271.38 ;
     RECT  349.06 305.2 350.3 317.58 ;
     RECT  349.34 381.22 350.5 698.98 ;
     RECT  349.82 255.22 350.98 271.38 ;
     RECT  346.66 146.44 351.94 165.96 ;
     RECT  350.3 304.36 351.94 317.58 ;
     RECT  343.1 335.44 351.94 354.96 ;
     RECT  346.94 205.24 352.9 236.94 ;
     RECT  347.9 283.36 352.9 292.38 ;
     RECT  350.5 386.68 352.9 698.98 ;
     RECT  351.94 342.58 353.18 354.96 ;
     RECT  353.18 342.58 353.38 361.68 ;
     RECT  352.9 283.36 355.3 289.44 ;
     RECT  352.9 226.24 356.06 236.94 ;
     RECT  352.9 386.68 356.26 415.06 ;
     RECT  351.94 305.2 357.7 316.74 ;
     RECT  356.06 226.24 357.98 237.36 ;
     RECT  357.7 305.2 358.66 309.6 ;
     RECT  356.26 386.68 359.14 391.92 ;
     RECT  350.98 259.84 359.62 271.38 ;
     RECT  357.98 226.24 361.06 240.3 ;
     RECT  359.14 391.72 361.54 391.92 ;
     RECT  353.38 343.42 362.02 361.68 ;
     RECT  356.54 251.02 362.5 251.22 ;
     RECT  356.54 280.42 362.5 280.62 ;
     RECT  362.02 361.48 362.98 361.68 ;
     RECT  356.26 401 362.98 415.06 ;
     RECT  355.3 289.24 363.26 289.44 ;
     RECT  351.94 146.44 363.46 161.76 ;
     RECT  363.26 289.24 364.42 294.9 ;
     RECT  352.9 205.24 364.9 214.26 ;
     RECT  359.62 264.46 364.9 271.38 ;
     RECT  364.9 271.18 366.14 271.38 ;
     RECT  362.78 322 366.82 322.2 ;
     RECT  358.66 308.56 367.1 309.6 ;
     RECT  365.66 248.5 367.3 248.7 ;
     RECT  361.06 226.24 367.78 239.46 ;
     RECT  366.14 271.18 367.78 272.64 ;
     RECT  364.9 205.24 368.06 205.44 ;
     RECT  367.1 307.72 368.06 309.6 ;
     RECT  367.1 318.64 368.06 318.84 ;
     RECT  368.06 198.1 368.26 205.44 ;
     RECT  367.78 227.5 368.26 239.46 ;
     RECT  367.78 271.18 368.26 271.38 ;
     RECT  364.42 289.24 368.26 289.44 ;
     RECT  362.02 343.42 368.26 352.02 ;
     RECT  368.06 307.72 368.74 318.84 ;
     RECT  364.9 214.06 369.22 214.26 ;
     RECT  362.98 401 369.5 414.64 ;
     RECT  368.26 349.3 370.46 352.02 ;
     RECT  369.02 385.84 370.46 386.04 ;
     RECT  369.5 168.28 370.94 168.48 ;
     RECT  368.54 337.12 371.62 339.84 ;
     RECT  370.46 349.3 372.1 358.32 ;
     RECT  352.9 424.1 372.58 698.98 ;
     RECT  369.5 400.54 372.86 414.64 ;
     RECT  368.06 369.04 373.06 369.24 ;
     RECT  372.58 428.3 373.06 652.78 ;
     RECT  363.46 146.44 373.34 154.2 ;
     RECT  368.74 307.72 373.34 316.74 ;
     RECT  373.06 428.3 373.54 651.52 ;
     RECT  370.94 168.28 373.82 169.32 ;
     RECT  368.06 258.16 373.82 258.36 ;
     RECT  368.54 124.18 374.02 124.38 ;
     RECT  373.82 165.76 374.02 169.32 ;
     RECT  373.34 146.44 374.3 156.72 ;
     RECT  372.38 285.04 374.78 285.24 ;
     RECT  372.1 349.72 375.26 358.32 ;
     RECT  374.02 165.76 375.46 168.9 ;
     RECT  371.62 339.64 375.46 339.84 ;
     RECT  372.86 188.44 375.74 188.64 ;
     RECT  374.3 146.44 376.22 157.14 ;
     RECT  371.42 113.26 376.7 113.46 ;
     RECT  373.82 258.16 377.18 267.18 ;
     RECT  373.34 305.62 377.18 316.74 ;
     RECT  375.74 184.66 377.66 188.64 ;
     RECT  375.26 349.72 378.34 362.1 ;
     RECT  377.18 305.62 378.62 320.1 ;
     RECT  368.26 227.5 379.58 227.7 ;
     RECT  368.26 239.26 379.58 239.46 ;
     RECT  374.78 283.78 379.58 285.24 ;
     RECT  376.7 112.84 379.78 113.46 ;
     RECT  370.46 385.84 380.06 391.08 ;
     RECT  372.86 399.7 380.06 414.64 ;
     RECT  377.18 258.16 380.74 269.7 ;
     RECT  379.58 283.78 381.02 286.08 ;
     RECT  377.66 180.88 381.7 188.64 ;
     RECT  379.58 239.26 381.7 241.14 ;
     RECT  381.7 240.94 382.18 241.14 ;
     RECT  373.54 433.76 382.94 651.52 ;
     RECT  372.58 662.66 382.94 698.98 ;
     RECT  378.62 305.62 383.14 327.24 ;
     RECT  375.74 127.12 383.9 127.32 ;
     RECT  376.22 138.88 383.9 157.14 ;
     RECT  382.94 433.76 384.86 698.98 ;
     RECT  383.9 127.12 385.06 157.14 ;
     RECT  381.02 283.78 385.34 286.92 ;
     RECT  385.06 130.9 385.82 157.14 ;
     RECT  375.46 165.76 385.82 166.8 ;
     RECT  380.06 385.84 386.3 414.64 ;
     RECT  378.34 354.34 387.46 362.1 ;
     RECT  386.3 379.96 387.74 414.64 ;
     RECT  381.7 188.44 388.7 188.64 ;
     RECT  368.26 198.1 388.7 205.02 ;
     RECT  385.82 130.9 389.18 166.8 ;
     RECT  379.58 222.46 389.18 227.7 ;
     RECT  385.34 283.78 390.14 287.76 ;
     RECT  385.34 297.64 390.14 298.68 ;
     RECT  388.7 188.44 391.58 205.02 ;
     RECT  389.18 222.46 391.58 230.22 ;
     RECT  383.14 308.98 391.58 327.24 ;
     RECT  389.18 130.9 391.78 172.68 ;
     RECT  390.14 283.78 392.54 298.68 ;
     RECT  391.58 307.3 392.54 327.24 ;
     RECT  387.74 377.02 392.74 414.64 ;
     RECT  379.78 112.84 393.22 113.04 ;
     RECT  392.54 283.78 393.22 327.24 ;
     RECT  391.58 222.04 393.98 230.22 ;
     RECT  391.58 182.14 394.94 205.02 ;
     RECT  391.78 130.9 395.14 168.48 ;
     RECT  392.74 377.02 396.1 407.88 ;
     RECT  394.94 182.14 396.58 211.74 ;
     RECT  380.74 258.16 396.86 267.6 ;
     RECT  396.86 258.16 397.06 275.16 ;
     RECT  393.98 222.04 397.34 235.26 ;
     RECT  386.3 101.5 398.98 101.7 ;
     RECT  384.86 427 399.26 698.98 ;
     RECT  397.06 258.16 399.46 274.74 ;
     RECT  397.34 222.04 400.22 241.14 ;
     RECT  395.14 130.9 400.42 158.4 ;
     RECT  397.34 340.48 400.9 340.68 ;
     RECT  396.1 392.56 400.9 407.88 ;
     RECT  400.22 222.04 402.14 244.92 ;
     RECT  399.26 422.8 402.14 698.98 ;
     RECT  402.14 222.04 402.62 247.02 ;
     RECT  400.9 392.56 402.82 403.68 ;
     RECT  402.14 422.38 403.1 698.98 ;
     RECT  402.62 222.04 403.3 248.28 ;
     RECT  399.46 258.16 403.3 267.6 ;
     RECT  403.3 235.06 403.78 248.28 ;
     RECT  393.22 283.78 404.54 287.34 ;
     RECT  393.22 297.64 404.54 327.24 ;
     RECT  396.1 377.02 404.54 381 ;
     RECT  395.14 168.28 405.22 168.48 ;
     RECT  404.54 283.78 405.7 327.24 ;
     RECT  403.1 418.6 405.7 698.98 ;
     RECT  396.58 196 406.66 211.74 ;
     RECT  405.7 283.78 407.14 286.08 ;
     RECT  402.82 394.66 407.62 403.68 ;
     RECT  403.3 222.04 408.1 222.24 ;
     RECT  407.14 283.78 408.1 285.24 ;
     RECT  406.66 199.36 408.58 211.74 ;
     RECT  405.7 299.74 408.58 327.24 ;
     RECT  408.58 206.92 408.86 211.74 ;
     RECT  403.3 267.4 408.86 267.6 ;
     RECT  408.86 267.4 409.54 272.64 ;
     RECT  408.86 206.92 410.02 218.04 ;
     RECT  408.58 301.84 410.02 327.24 ;
     RECT  409.54 272.44 410.5 272.64 ;
     RECT  400.42 146.44 410.98 158.4 ;
     RECT  403.78 235.06 411.46 247.44 ;
     RECT  408.1 285.04 412.42 285.24 ;
     RECT  410.02 206.92 412.9 207.12 ;
     RECT  411.46 244.72 413.86 247.44 ;
     RECT  403.3 258.16 413.86 258.36 ;
     RECT  407.62 396.76 413.86 403.68 ;
     RECT  404.54 377.02 414.14 381.42 ;
     RECT  400.42 130.9 414.82 131.1 ;
     RECT  414.14 377.02 415.3 383.1 ;
     RECT  411.74 172.9 415.78 173.1 ;
     RECT  415.3 379.96 415.78 383.1 ;
     RECT  411.46 235.06 416.06 235.26 ;
     RECT  410.98 146.44 416.26 156.72 ;
     RECT  416.06 232.54 416.26 235.26 ;
     RECT  410.02 301.84 416.26 325.14 ;
     RECT  416.26 301.84 416.74 302.04 ;
     RECT  416.26 156.52 417.22 156.72 ;
     RECT  413.86 244.72 417.22 244.92 ;
     RECT  416.26 146.44 417.98 147.06 ;
     RECT  396.58 182.14 417.98 182.34 ;
     RECT  413.66 347.2 417.98 347.4 ;
     RECT  410.02 217.84 418.18 218.04 ;
     RECT  413.86 397.6 418.18 403.68 ;
     RECT  417.98 175 418.46 182.34 ;
     RECT  417.98 343 418.46 348.66 ;
     RECT  416.26 232.54 418.66 232.74 ;
     RECT  418.46 343 418.94 349.08 ;
     RECT  410.78 366.94 418.94 367.14 ;
     RECT  418.46 175 419.62 184.86 ;
     RECT  419.42 287.56 419.9 288.18 ;
     RECT  418.94 365.68 419.9 367.14 ;
     RECT  419.62 180.88 420.1 182.76 ;
     RECT  418.94 343 420.38 349.5 ;
     RECT  419.9 360.64 420.38 367.14 ;
     RECT  420.38 343 420.86 367.14 ;
     RECT  419.9 287.56 421.82 288.6 ;
     RECT  420.86 337.96 422.02 367.14 ;
     RECT  422.02 338.8 422.3 367.14 ;
     RECT  421.82 285.04 422.78 288.6 ;
     RECT  421.34 297.22 422.78 297.42 ;
     RECT  418.18 397.6 422.78 397.8 ;
     RECT  423.26 266.98 423.74 267.18 ;
     RECT  422.78 285.04 424.22 297.42 ;
     RECT  421.34 407.26 424.22 407.46 ;
     RECT  405.7 422.38 424.22 698.98 ;
     RECT  422.78 395.08 424.42 397.8 ;
     RECT  422.3 228.34 426.34 228.54 ;
     RECT  424.22 279.16 426.34 297.42 ;
     RECT  422.3 338.8 426.34 367.98 ;
     RECT  423.26 123.76 426.82 123.96 ;
     RECT  416.26 310.66 427.1 325.14 ;
     RECT  417.98 142.66 427.3 147.06 ;
     RECT  415.78 379.96 427.78 380.16 ;
     RECT  420.38 162.4 428.06 162.6 ;
     RECT  423.74 259.84 428.06 267.18 ;
     RECT  427.1 308.98 428.26 325.14 ;
     RECT  428.06 259.84 428.74 275.58 ;
     RECT  419.9 211.12 429.02 211.32 ;
     RECT  424.22 407.26 429.02 698.98 ;
     RECT  429.02 399.7 429.22 698.98 ;
     RECT  428.06 161.56 429.5 162.6 ;
     RECT  429.02 207.34 429.5 211.32 ;
     RECT  429.5 207.34 429.98 214.68 ;
     RECT  428.26 310.66 429.98 325.14 ;
     RECT  426.34 338.8 430.18 365.88 ;
     RECT  429.98 310.66 431.14 328.92 ;
     RECT  427.3 142.66 431.62 146.64 ;
     RECT  426.34 284.2 431.9 297.42 ;
     RECT  431.62 143.5 432.1 146.64 ;
     RECT  431.14 310.66 432.1 325.14 ;
     RECT  430.18 339.22 432.1 365.88 ;
     RECT  429.5 161.56 432.58 166.8 ;
     RECT  420.1 180.88 432.58 182.34 ;
     RECT  428.74 266.98 433.06 275.58 ;
     RECT  429.98 207.34 433.82 215.1 ;
     RECT  431.9 284.2 435.94 299.1 ;
     RECT  418.46 100.66 436.9 100.86 ;
     RECT  432.1 310.66 436.9 320.94 ;
     RECT  435.94 284.2 437.38 294.06 ;
     RECT  438.14 249.76 439.1 249.96 ;
     RECT  433.82 206.08 439.3 215.1 ;
     RECT  432.1 339.22 439.3 362.94 ;
     RECT  433.06 266.98 439.78 271.38 ;
     RECT  439.3 206.08 440.26 211.32 ;
     RECT  439.1 127.54 440.54 127.74 ;
     RECT  432.1 146.44 441.5 146.64 ;
     RECT  440.54 373.66 441.5 373.86 ;
     RECT  432.58 162.4 441.7 166.8 ;
     RECT  429.22 415.66 442.18 698.98 ;
     RECT  439.1 249.76 442.46 253.74 ;
     RECT  439.78 271.18 442.46 271.38 ;
     RECT  437.38 284.2 442.46 288.18 ;
     RECT  439.3 339.22 442.46 362.52 ;
     RECT  429.22 399.7 443.14 399.9 ;
     RECT  436.7 225.82 443.42 226.02 ;
     RECT  441.5 373.24 443.62 373.86 ;
     RECT  442.46 246.82 446.3 253.74 ;
     RECT  442.46 271.18 446.98 288.18 ;
     RECT  442.18 422.38 447.46 698.98 ;
     RECT  446.98 284.2 447.74 288.18 ;
     RECT  443.42 225.82 449.18 232.32 ;
     RECT  446.3 246.82 449.18 254.16 ;
     RECT  442.46 338.8 449.86 362.52 ;
     RECT  436.9 312.76 450.14 320.52 ;
     RECT  432.58 182.14 450.34 182.34 ;
     RECT  450.14 312.76 450.34 327.66 ;
     RECT  441.5 138.88 451.78 146.64 ;
     RECT  450.34 314.44 451.78 327.66 ;
     RECT  449.86 345.94 451.78 362.52 ;
     RECT  440.54 120.82 452.74 127.74 ;
     RECT  451.78 146.44 453.22 146.64 ;
     RECT  451.78 314.44 453.22 322.62 ;
     RECT  447.74 284.2 453.98 290.28 ;
     RECT  453.22 314.86 454.18 322.62 ;
     RECT  451.78 348.88 454.18 362.52 ;
     RECT  454.18 348.88 454.66 357.48 ;
     RECT  449.18 225.82 454.94 254.16 ;
     RECT  453.98 284.2 454.94 296.58 ;
     RECT  442.94 388.78 454.94 388.98 ;
     RECT  454.94 225.82 455.14 259.62 ;
     RECT  454.66 350.14 455.14 357.48 ;
     RECT  455.14 245.56 455.62 259.62 ;
     RECT  455.62 245.98 456.1 259.62 ;
     RECT  455.14 225.82 456.58 232.32 ;
     RECT  447.46 422.38 459.26 587.68 ;
     RECT  447.46 597.56 459.26 698.98 ;
     RECT  454.94 284.2 460.42 298.26 ;
     RECT  460.42 284.2 460.9 296.16 ;
     RECT  452.74 120.82 461.38 121.02 ;
     RECT  456.58 225.82 461.38 226.02 ;
     RECT  454.18 314.86 463.1 320.1 ;
     RECT  456.1 248.92 463.3 259.62 ;
     RECT  443.62 373.66 463.3 373.86 ;
     RECT  459.26 422.38 463.3 698.98 ;
     RECT  463.3 257.32 463.78 259.62 ;
     RECT  460.9 284.2 463.78 290.28 ;
     RECT  441.7 166.6 465.22 166.8 ;
     RECT  454.94 383.74 465.22 388.98 ;
     RECT  463.1 306.46 465.5 320.1 ;
     RECT  464.54 282.94 466.18 283.56 ;
     RECT  465.5 306.46 466.66 325.14 ;
     RECT  465.22 384.58 466.66 388.98 ;
     RECT  440.26 211.12 467.14 211.32 ;
     RECT  455.14 350.14 467.62 350.34 ;
     RECT  457.82 154.84 468.1 155.04 ;
     RECT  463.78 257.32 468.1 257.52 ;
     RECT  466.66 306.46 468.86 320.94 ;
     RECT  464.54 248.5 469.06 248.7 ;
     RECT  465.02 369.46 469.06 369.66 ;
     RECT  463.3 422.38 469.54 653.2 ;
     RECT  469.54 576.14 470.02 653.2 ;
     RECT  468.86 212.8 471.26 220.98 ;
     RECT  469.34 332.5 471.74 333.54 ;
     RECT  468.86 282.52 472.22 282.72 ;
     RECT  470.02 580.76 472.7 653.2 ;
     RECT  463.3 662.66 472.7 698.98 ;
     RECT  472.22 279.58 474.14 282.72 ;
     RECT  470.78 181.3 474.34 181.5 ;
     RECT  471.74 162.4 475.3 162.6 ;
     RECT  468.86 301 475.3 320.94 ;
     RECT  475.3 301.42 476.26 320.94 ;
     RECT  474.14 279.16 477.02 282.72 ;
     RECT  476.06 195.58 477.5 195.78 ;
     RECT  477.5 377.44 477.98 377.64 ;
     RECT  471.74 332.5 478.46 337.32 ;
     RECT  470.78 347.2 478.46 347.4 ;
     RECT  474.62 241.36 479.42 241.56 ;
     RECT  478.46 332.5 479.42 347.4 ;
     RECT  472.7 116.2 479.62 116.4 ;
     RECT  479.42 241.36 479.9 241.98 ;
     RECT  477.02 277.06 480.38 282.72 ;
     RECT  477.5 188.02 481.06 195.78 ;
     RECT  480.38 272.44 482.02 282.72 ;
     RECT  479.9 241.36 482.78 244.92 ;
     RECT  478.46 256.06 482.78 256.26 ;
     RECT  476.26 304.36 482.78 320.94 ;
     RECT  479.42 332.5 482.78 354.96 ;
     RECT  482.78 241.36 482.98 256.26 ;
     RECT  476.54 130.06 484.42 130.26 ;
     RECT  482.78 177.1 484.42 177.3 ;
     RECT  482.78 304.36 484.42 354.96 ;
     RECT  471.26 212.8 485.18 223.08 ;
     RECT  482.02 277.06 486.62 282.72 ;
     RECT  483.74 294.7 486.62 294.9 ;
     RECT  479.9 368.62 487.58 368.82 ;
     RECT  477.98 377.44 487.58 385.2 ;
     RECT  469.54 422.38 488.74 565.84 ;
     RECT  485.18 212.8 489.5 226.86 ;
     RECT  482.98 241.36 489.5 248.7 ;
     RECT  489.5 212.8 490.66 248.7 ;
     RECT  472.7 580.76 490.66 698.98 ;
     RECT  483.74 263.2 492.1 263.4 ;
     RECT  488.74 422.38 493.54 545.26 ;
     RECT  491.42 131.32 493.82 131.52 ;
     RECT  484.42 308.56 493.82 354.96 ;
     RECT  493.82 131.32 494.02 132.36 ;
     RECT  490.66 241.36 494.02 248.7 ;
     RECT  494.02 131.32 494.78 131.94 ;
     RECT  494.02 241.78 494.98 248.7 ;
     RECT  478.94 161.56 495.26 161.76 ;
     RECT  486.62 277.06 495.26 294.9 ;
     RECT  493.82 304.36 495.26 354.96 ;
     RECT  495.26 161.56 495.46 169.74 ;
     RECT  481.06 195.58 495.46 195.78 ;
     RECT  494.98 248.5 495.74 248.7 ;
     RECT  495.26 277.06 496.42 354.96 ;
     RECT  493.54 422.38 497.38 537.7 ;
     RECT  490.66 212.8 498.14 229.8 ;
     RECT  498.14 204.82 498.34 229.8 ;
     RECT  496.42 277.06 498.82 304.98 ;
     RECT  494.78 130.9 499.78 131.94 ;
     RECT  498.82 300.58 501.22 304.98 ;
     RECT  487.58 368.62 501.22 388.98 ;
     RECT  501.22 301.84 501.7 304.98 ;
     RECT  493.34 109.06 502.18 109.26 ;
     RECT  493.82 185.08 502.94 185.28 ;
     RECT  498.34 220.78 503.42 229.8 ;
     RECT  490.66 588.32 503.62 698.98 ;
     RECT  492.86 399.7 505.06 399.9 ;
     RECT  495.74 248.5 505.34 251.22 ;
     RECT  503.62 588.32 505.34 652.36 ;
     RECT  502.94 180.88 505.54 185.28 ;
     RECT  497.38 422.38 505.54 425.1 ;
     RECT  505.34 583.7 506.02 652.36 ;
     RECT  495.46 167.86 506.5 169.74 ;
     RECT  503.42 220.78 506.5 232.74 ;
     RECT  488.74 557.24 506.78 565.84 ;
     RECT  498.34 204.82 506.98 205.02 ;
     RECT  503.62 662.24 506.98 698.98 ;
     RECT  506.5 169.54 507.46 169.74 ;
     RECT  505.34 248.5 507.46 253.74 ;
     RECT  496.42 314.86 507.94 354.96 ;
     RECT  506.78 555.56 508.22 565.84 ;
     RECT  506.78 120.4 509.38 120.6 ;
     RECT  506.5 222.46 509.38 232.74 ;
     RECT  505.54 422.38 509.86 422.58 ;
     RECT  507.46 248.5 511.3 248.7 ;
     RECT  499.78 130.9 512.06 131.52 ;
     RECT  498.82 277.06 512.54 290.7 ;
     RECT  507.94 314.86 512.54 351.18 ;
     RECT  512.54 276.64 513.02 290.7 ;
     RECT  512.06 130.9 513.22 135.3 ;
     RECT  506.02 583.7 513.5 646.06 ;
     RECT  513.02 272.44 514.18 290.7 ;
     RECT  501.22 369.46 514.46 388.98 ;
     RECT  508.22 555.56 514.46 568.36 ;
     RECT  513.5 577.4 514.46 646.06 ;
     RECT  501.7 301.84 514.94 302.04 ;
     RECT  512.54 312.76 514.94 351.18 ;
     RECT  514.46 555.56 514.94 646.06 ;
     RECT  509.38 222.46 515.14 222.66 ;
     RECT  514.94 301.84 515.14 351.18 ;
     RECT  497.38 433.76 515.14 537.7 ;
     RECT  514.46 369.04 516.1 390.66 ;
     RECT  514.18 276.64 516.38 290.7 ;
     RECT  515.14 301.84 516.38 344.88 ;
     RECT  510.62 116.2 516.58 116.4 ;
     RECT  514.94 549.26 516.58 646.06 ;
     RECT  516.1 369.04 516.86 390.24 ;
     RECT  506.98 662.66 516.86 698.98 ;
     RECT  516.86 366.1 517.54 390.24 ;
     RECT  505.54 180.88 518.02 181.08 ;
     RECT  516.38 276.64 518.02 344.88 ;
     RECT  513.22 135.1 518.5 135.3 ;
     RECT  518.02 276.64 518.5 283.14 ;
     RECT  516.58 549.26 518.5 592.72 ;
     RECT  517.54 383.74 518.98 390.24 ;
     RECT  505.82 154.42 519.26 154.62 ;
     RECT  509.38 232.54 519.26 232.74 ;
     RECT  511.58 241.78 519.46 241.98 ;
     RECT  518.02 297.22 519.46 344.88 ;
     RECT  519.26 232.54 519.74 233.16 ;
     RECT  519.74 232.54 520.22 234 ;
     RECT  516.86 407.26 520.7 407.46 ;
     RECT  518.5 549.26 520.7 591.88 ;
     RECT  519.26 146.02 521.66 154.62 ;
     RECT  520.7 165.76 521.66 165.96 ;
     RECT  521.18 206.08 522.34 210.48 ;
     RECT  516.58 632 522.34 646.06 ;
     RECT  519.46 298.06 523.78 304.56 ;
     RECT  521.66 146.02 524.54 165.96 ;
     RECT  518.5 276.64 524.54 278.94 ;
     RECT  523.78 304.36 525.22 304.56 ;
     RECT  522.34 632 525.5 645.64 ;
     RECT  517.54 366.1 525.7 369.66 ;
     RECT  524.54 146.02 526.18 170.16 ;
     RECT  524.54 272.44 526.18 278.94 ;
     RECT  516.58 602.18 526.18 622.96 ;
     RECT  524.54 188.02 526.46 188.22 ;
     RECT  520.22 229.6 526.94 234 ;
     RECT  525.7 369.46 526.94 369.66 ;
     RECT  520.7 547.16 526.94 591.88 ;
     RECT  526.18 276.64 527.14 278.94 ;
     RECT  526.94 369.46 527.62 373.44 ;
     RECT  522.34 206.08 528.1 206.28 ;
     RECT  515.14 433.76 528.86 536.44 ;
     RECT  526.94 545.48 528.86 591.88 ;
     RECT  520.7 399.7 529.54 407.46 ;
     RECT  527.42 279.16 529.82 279.36 ;
     RECT  528.86 433.76 530.3 591.88 ;
     RECT  523.1 119.98 531.46 120.18 ;
     RECT  525.5 631.58 531.46 645.64 ;
     RECT  530.3 305.2 531.74 305.4 ;
     RECT  519.46 317.38 531.74 332.28 ;
     RECT  521.66 354.76 531.74 354.96 ;
     RECT  526.94 222.04 532.22 234 ;
     RECT  522.62 131.74 532.7 131.94 ;
     RECT  516.86 655.52 532.9 698.98 ;
     RECT  532.22 222.04 533.38 238.62 ;
     RECT  532.7 131.74 533.66 135.3 ;
     RECT  527.62 372.82 534.14 373.44 ;
     RECT  518.98 383.74 534.14 383.94 ;
     RECT  530.3 433.76 534.14 593.14 ;
     RECT  526.18 602.18 534.14 618.34 ;
     RECT  531.46 632 534.34 645.64 ;
     RECT  526.46 180.88 534.82 188.22 ;
     RECT  531.74 354.34 534.82 354.96 ;
     RECT  526.18 150.22 535.3 170.16 ;
     RECT  531.74 305.2 536.26 332.28 ;
     RECT  534.14 372.82 536.74 388.98 ;
     RECT  536.26 319.9 537.02 332.28 ;
     RECT  519.46 342.16 537.02 344.88 ;
     RECT  536.74 387.94 537.02 388.98 ;
     RECT  535.3 158.2 537.7 170.16 ;
     RECT  533.66 131.74 538.46 135.72 ;
     RECT  534.14 433.76 539.14 618.34 ;
     RECT  537.7 158.2 539.62 165.96 ;
     RECT  538.46 131.74 540.38 143.28 ;
     RECT  537.02 319.9 540.38 344.88 ;
     RECT  534.82 354.34 540.38 354.54 ;
     RECT  539.14 434.6 540.58 618.34 ;
     RECT  529.82 279.16 541.34 283.98 ;
     RECT  533.38 222.04 541.54 230.64 ;
     RECT  541.34 279.16 541.54 290.7 ;
     RECT  529.54 407.26 541.54 407.46 ;
     RECT  534.82 188.02 542.98 188.22 ;
     RECT  538.94 268.24 542.98 268.44 ;
     RECT  532.9 662.66 542.98 698.98 ;
     RECT  540.58 435.44 543.46 618.34 ;
     RECT  534.34 632 543.46 645.22 ;
     RECT  537.02 387.94 544.42 392.34 ;
     RECT  540.38 131.32 544.7 143.28 ;
     RECT  536.74 372.82 545.18 373.02 ;
     RECT  539.62 165.76 546.34 165.96 ;
     RECT  536.26 305.2 546.34 309.18 ;
     RECT  540.38 319.9 546.34 354.54 ;
     RECT  543.46 435.44 546.34 614.98 ;
     RECT  542.78 199.78 546.62 199.98 ;
     RECT  537.5 105.28 547.3 105.48 ;
     RECT  546.62 199.78 548.06 203.76 ;
     RECT  544.42 392.14 549.22 392.34 ;
     RECT  532.7 248.92 549.98 249.12 ;
     RECT  549.02 260.26 549.98 260.46 ;
     RECT  546.34 347.2 549.98 354.54 ;
     RECT  545.18 372.82 549.98 376.8 ;
     RECT  546.34 319.9 550.46 331.86 ;
     RECT  546.34 441.32 550.66 614.98 ;
     RECT  541.54 279.16 551.14 279.36 ;
     RECT  549.98 347.2 551.62 357.06 ;
     RECT  549.98 372.82 551.62 377.64 ;
     RECT  546.34 305.2 552.58 305.4 ;
     RECT  542.98 662.66 552.58 697.72 ;
     RECT  549.98 248.92 553.06 260.46 ;
     RECT  544.7 131.32 553.34 146.64 ;
     RECT  553.06 248.92 553.54 249.12 ;
     RECT  550.66 444.26 554.5 614.98 ;
     RECT  543.46 644.18 554.5 645.22 ;
     RECT  550.46 316.54 555.46 331.86 ;
     RECT  551.62 347.2 555.46 354.54 ;
     RECT  549.02 161.98 557.18 162.18 ;
     RECT  553.34 122.92 557.38 146.64 ;
     RECT  548.06 199.78 557.66 207.54 ;
     RECT  557.38 122.92 557.86 131.94 ;
     RECT  557.66 196 557.86 207.54 ;
     RECT  553.06 260.26 558.82 260.46 ;
     RECT  554.5 454.76 558.82 614.98 ;
     RECT  541.54 222.04 559.58 222.24 ;
     RECT  551.9 233.38 559.58 233.58 ;
     RECT  555.46 354.34 559.78 354.54 ;
     RECT  557.18 161.98 562.18 165.96 ;
     RECT  559.58 222.04 562.18 233.58 ;
     RECT  557.38 143.08 562.66 146.64 ;
     RECT  557.86 196 562.94 199.56 ;
     RECT  554.78 273.7 562.94 274.32 ;
     RECT  562.94 194.74 563.14 199.56 ;
     RECT  562.18 161.98 564.1 162.18 ;
     RECT  554.5 644.18 564.1 644.8 ;
     RECT  557.86 122.92 564.58 123.96 ;
     RECT  562.66 143.08 565.06 143.28 ;
     RECT  562.18 227.08 565.06 233.58 ;
     RECT  562.94 273.7 565.34 281.88 ;
     RECT  541.54 290.5 565.34 290.7 ;
     RECT  564.58 123.76 566.5 123.96 ;
     RECT  565.34 273.7 566.5 290.7 ;
     RECT  566.5 273.7 566.98 278.1 ;
     RECT  563.14 196 568.42 199.56 ;
     RECT  566.78 300.16 568.9 300.36 ;
     RECT  555.46 316.54 569.66 328.92 ;
     RECT  554.5 444.26 569.66 445.72 ;
     RECT  558.82 454.76 569.66 614.14 ;
     RECT  569.66 308.98 569.86 330.6 ;
     RECT  569.86 320.32 570.82 320.94 ;
     RECT  552.58 662.66 572.06 696.88 ;
     RECT  568.22 247.66 573.98 247.86 ;
     RECT  564.1 644.18 573.98 644.38 ;
     RECT  565.06 227.08 575.62 229.38 ;
     RECT  573.98 241.36 575.62 247.86 ;
     RECT  569.66 444.26 576.1 614.14 ;
     RECT  571.1 173.32 576.38 173.52 ;
     RECT  576.1 444.26 577.06 445.72 ;
     RECT  576.38 169.12 577.34 173.52 ;
     RECT  570.14 199.78 577.34 199.98 ;
     RECT  570.62 297.64 577.34 297.84 ;
     RECT  569.86 308.98 577.34 309.18 ;
     RECT  575.62 229.18 577.54 229.38 ;
     RECT  574.46 339.22 577.54 345.72 ;
     RECT  570.62 622.76 577.82 622.96 ;
     RECT  543.46 632 577.82 632.2 ;
     RECT  567.26 135.52 578.3 138.66 ;
     RECT  566.98 274.54 578.3 278.1 ;
     RECT  569.86 330.4 578.3 330.6 ;
     RECT  577.54 339.22 578.3 339.42 ;
     RECT  569.66 379.96 578.3 380.16 ;
     RECT  576.86 388.78 578.3 388.98 ;
     RECT  578.3 131.32 578.5 138.66 ;
     RECT  577.34 199.78 578.5 201.66 ;
     RECT  571.58 154.42 579.26 154.62 ;
     RECT  577.34 169.12 579.26 178.56 ;
     RECT  577.82 622.76 579.26 633.04 ;
     RECT  573.98 643.76 579.26 644.38 ;
     RECT  572.06 654.26 579.46 696.88 ;
     RECT  575.42 358.12 580.22 358.32 ;
     RECT  570.82 320.32 580.42 320.52 ;
     RECT  580.22 350.56 580.42 358.32 ;
     RECT  578.3 379.96 580.9 388.98 ;
     RECT  576.1 456.02 581.38 614.14 ;
     RECT  579.26 168.7 581.66 178.56 ;
     RECT  577.34 297.64 583.1 309.18 ;
     RECT  583.1 297.64 584.54 313.38 ;
     RECT  577.06 445.52 584.74 445.72 ;
     RECT  581.38 456.02 584.74 607 ;
     RECT  575.62 247.66 585.22 247.86 ;
     RECT  584.74 456.02 585.22 603.64 ;
     RECT  578.5 199.78 585.5 199.98 ;
     RECT  585.22 544.64 585.7 603.64 ;
     RECT  578.3 274.54 586.94 278.94 ;
     RECT  584.54 291.34 587.14 313.38 ;
     RECT  580.42 350.56 587.62 351.18 ;
     RECT  585.7 546.32 587.62 603.64 ;
     RECT  579.74 230.02 587.9 234 ;
     RECT  586.94 274.54 587.9 282.3 ;
     RECT  585.5 196 588.1 199.98 ;
     RECT  579.26 622.76 588.38 644.38 ;
     RECT  588.1 199.78 588.58 199.98 ;
     RECT  587.14 294.28 588.58 313.38 ;
     RECT  585.22 456.02 589.54 535.18 ;
     RECT  587.9 230.02 589.82 237.36 ;
     RECT  589.54 456.02 590.02 502.42 ;
     RECT  578.3 330.4 590.3 339.42 ;
     RECT  587.62 350.56 590.3 350.76 ;
     RECT  578.5 131.32 590.5 136.14 ;
     RECT  587.62 551.78 590.5 603.64 ;
     RECT  579.26 153.16 591.26 154.62 ;
     RECT  581.66 168.28 591.26 178.56 ;
     RECT  591.26 153.16 591.46 178.56 ;
     RECT  585.5 369.88 592.7 370.08 ;
     RECT  590.5 131.32 592.9 135.72 ;
     RECT  588.86 264.04 594.14 264.24 ;
     RECT  587.9 274.12 594.14 282.3 ;
     RECT  590.3 330.4 594.14 350.76 ;
     RECT  589.82 226.24 595.3 237.36 ;
     RECT  580.9 379.96 595.3 385.2 ;
     RECT  590.02 456.02 595.3 500.74 ;
     RECT  595.3 230.02 595.78 237.36 ;
     RECT  588.38 617.72 595.78 644.38 ;
     RECT  592.7 366.1 596.06 370.08 ;
     RECT  595.3 379.96 596.06 381.42 ;
     RECT  595.78 230.02 596.26 234.42 ;
     RECT  595.3 468.62 596.26 500.74 ;
     RECT  591.46 161.98 596.74 178.56 ;
     RECT  595.3 456.02 596.74 456.22 ;
     RECT  579.46 655.94 596.74 696.88 ;
     RECT  588.58 297.64 597.22 313.38 ;
     RECT  595.78 621.08 597.22 644.38 ;
     RECT  597.22 313.18 597.7 313.38 ;
     RECT  590.5 551.78 597.7 590.2 ;
     RECT  593.66 252.7 598.66 252.9 ;
     RECT  597.7 577.82 598.66 590.2 ;
     RECT  596.26 468.62 599.14 483.1 ;
     RECT  598.66 583.7 599.14 590.2 ;
     RECT  590.5 598.82 599.14 603.64 ;
     RECT  588.86 395.92 599.42 396.12 ;
     RECT  592.9 131.74 599.62 135.72 ;
     RECT  596.26 491.72 599.62 500.74 ;
     RECT  599.14 481.22 600.1 483.1 ;
     RECT  597.98 192.22 600.58 196.62 ;
     RECT  599.14 468.62 601.06 472.6 ;
     RECT  597.22 632 601.06 644.38 ;
     RECT  594.14 264.04 601.34 282.3 ;
     RECT  601.34 264.04 601.54 286.5 ;
     RECT  597.22 621.08 601.54 622.96 ;
     RECT  597.02 207.34 602.02 207.54 ;
     RECT  600.1 482.06 602.02 483.1 ;
     RECT  594.14 327.88 602.3 350.76 ;
     RECT  599.62 491.72 602.5 496.96 ;
     RECT  599.14 583.7 602.5 583.9 ;
     RECT  589.54 515.24 602.98 535.18 ;
     RECT  601.06 470.3 603.46 470.5 ;
     RECT  602.02 482.48 603.46 483.1 ;
     RECT  596.74 662.66 603.46 696.88 ;
     RECT  603.46 482.48 604.42 482.68 ;
     RECT  600.58 192.22 604.9 192.42 ;
     RECT  602.3 327.88 605.38 354.54 ;
     RECT  605.38 327.88 605.86 342.36 ;
     RECT  599.42 395.92 606.14 396.54 ;
     RECT  597.22 297.64 606.34 301.62 ;
     RECT  596.06 366.1 606.34 381.42 ;
     RECT  599.14 598.82 606.34 599.02 ;
     RECT  601.54 269.08 606.82 286.5 ;
     RECT  591.46 153.16 607.3 153.36 ;
     RECT  602.98 515.24 607.3 530.56 ;
     RECT  601.54 621.08 608.06 621.28 ;
     RECT  606.14 395.92 608.26 402 ;
     RECT  605.66 312.34 608.54 312.54 ;
     RECT  608.06 613.52 609.22 621.28 ;
     RECT  596.74 162.4 609.5 178.56 ;
     RECT  606.34 300.16 609.7 301.62 ;
     RECT  608.54 312.34 610.18 316.32 ;
     RECT  606.34 369.88 610.18 381.42 ;
     RECT  603.46 663.08 610.66 696.88 ;
     RECT  597.7 551.78 611.42 565.84 ;
     RECT  611.42 252.7 611.62 253.32 ;
     RECT  611.42 545.9 611.62 565.84 ;
     RECT  596.26 230.02 612.1 234 ;
     RECT  611.62 565.64 612.38 565.84 ;
     RECT  609.7 300.16 612.58 300.36 ;
     RECT  608.26 395.92 612.58 396.54 ;
     RECT  601.06 632 612.86 632.2 ;
     RECT  610.18 369.88 613.06 375.96 ;
     RECT  601.06 644.18 613.34 644.38 ;
     RECT  609.5 160.72 613.54 178.56 ;
     RECT  599.62 132.58 614.3 135.72 ;
     RECT  612.1 233.8 614.98 234 ;
     RECT  613.34 644.18 615.46 644.8 ;
     RECT  612.86 630.74 615.74 632.2 ;
     RECT  613.54 160.72 615.94 160.92 ;
     RECT  606.82 269.08 615.94 282.3 ;
     RECT  610.18 316.12 615.94 316.32 ;
     RECT  605.86 327.88 616.7 337.74 ;
     RECT  614.3 131.74 616.9 139.5 ;
     RECT  612.58 396.34 617.38 396.54 ;
     RECT  612.38 565.64 617.38 569.2 ;
     RECT  611.62 545.9 618.14 551.98 ;
     RECT  616.9 131.74 618.34 131.94 ;
     RECT  613.06 369.88 618.82 374.28 ;
     RECT  611.9 595.46 619.1 595.66 ;
     RECT  611.62 253.12 619.58 253.32 ;
     RECT  615.94 272.02 619.78 282.3 ;
     RECT  619.78 274.12 620.06 282.3 ;
     RECT  619.1 595.46 620.06 596.08 ;
     RECT  620.06 274.12 620.26 282.72 ;
     RECT  616.7 324.1 620.26 337.74 ;
     RECT  615.74 630.74 620.54 633.04 ;
     RECT  620.06 197.26 622.18 197.46 ;
     RECT  619.58 253.12 622.18 256.26 ;
     RECT  609.22 613.52 622.18 613.72 ;
     RECT  617.38 565.64 622.46 566.26 ;
     RECT  620.54 626.96 622.66 633.04 ;
     RECT  613.54 172.9 622.94 178.56 ;
     RECT  618.82 373.24 622.94 374.28 ;
     RECT  620.54 383.74 622.94 383.94 ;
     RECT  610.66 666.86 624.58 696.88 ;
     RECT  621.5 240.94 624.86 241.14 ;
     RECT  621.02 146.86 625.34 147.06 ;
     RECT  605.38 354.34 625.34 354.54 ;
     RECT  624.86 240.94 626.02 248.28 ;
     RECT  618.14 545.48 626.02 551.98 ;
     RECT  625.34 146.86 626.3 147.48 ;
     RECT  623.42 158.2 626.3 158.4 ;
     RECT  622.94 172.9 626.3 188.64 ;
     RECT  624.38 313.18 626.3 313.38 ;
     RECT  620.26 324.1 626.3 333.96 ;
     RECT  620.06 294.28 626.78 297 ;
     RECT  625.34 349.72 626.78 354.54 ;
     RECT  626.78 349.72 627.26 354.96 ;
     RECT  626.3 146.86 627.46 158.4 ;
     RECT  627.26 349.72 627.74 358.74 ;
     RECT  620.06 595.04 627.94 596.08 ;
     RECT  623.42 131.32 628.22 131.52 ;
     RECT  626.78 294.28 628.22 301.2 ;
     RECT  626.3 313.18 628.22 333.96 ;
     RECT  627.46 146.86 628.9 154.62 ;
     RECT  623.42 203.14 628.9 203.34 ;
     RECT  626.02 240.94 629.18 244.92 ;
     RECT  620.26 282.52 629.18 282.72 ;
     RECT  628.22 291.34 629.18 333.96 ;
     RECT  622.94 373.24 629.18 383.94 ;
     RECT  629.18 291.34 629.86 340.26 ;
     RECT  609.5 584.12 629.86 584.32 ;
     RECT  629.86 316.96 630.14 340.26 ;
     RECT  627.74 349.72 630.14 359.58 ;
     RECT  629.18 370.3 630.34 383.94 ;
     RECT  622.46 564.8 630.34 566.26 ;
     RECT  629.18 278.74 630.62 282.72 ;
     RECT  629.86 291.34 630.82 305.82 ;
     RECT  625.82 264.04 631.1 264.24 ;
     RECT  627.94 595.04 631.1 595.66 ;
     RECT  602.5 491.72 631.3 494.44 ;
     RECT  630.62 275.38 631.58 282.72 ;
     RECT  630.82 291.34 631.58 301.2 ;
     RECT  630.14 316.96 631.58 359.58 ;
     RECT  626.3 170.38 631.78 188.64 ;
     RECT  629.18 236.32 631.78 244.92 ;
     RECT  631.78 172.9 632.74 188.64 ;
     RECT  631.58 275.38 632.74 301.2 ;
     RECT  631.1 587.9 632.74 595.66 ;
     RECT  628.9 153.58 633.22 154.62 ;
     RECT  623.42 607.22 633.7 607.42 ;
     RECT  615.46 644.18 633.98 644.38 ;
     RECT  631.78 237.16 634.18 244.92 ;
     RECT  632.74 595.46 634.18 595.66 ;
     RECT  632.74 172.9 635.14 184.86 ;
     RECT  632.74 296.8 635.14 301.2 ;
     RECT  607.3 515.24 635.14 529.3 ;
     RECT  633.22 153.58 635.62 153.78 ;
     RECT  635.14 172.9 635.62 176.88 ;
     RECT  631.58 316.96 635.9 361.68 ;
     RECT  630.34 370.3 635.9 378.06 ;
     RECT  628.22 131.32 636.1 135.72 ;
     RECT  635.9 316.96 636.58 378.06 ;
     RECT  626.02 545.48 636.58 550.3 ;
     RECT  636.58 316.96 637.06 340.26 ;
     RECT  636.1 135.52 637.54 135.72 ;
     RECT  635.14 301 637.54 301.2 ;
     RECT  637.06 316.96 637.54 335.64 ;
     RECT  634.18 244.72 638.5 244.92 ;
     RECT  631.3 491.72 638.5 491.92 ;
     RECT  633.98 644.18 638.5 652.78 ;
     RECT  631.1 260.26 638.78 264.24 ;
     RECT  636.58 550.1 640.42 550.3 ;
     RECT  622.66 632.84 641.38 633.04 ;
     RECT  637.54 316.96 641.66 317.16 ;
     RECT  637.54 327.88 641.86 335.64 ;
     RECT  636.58 349.72 641.86 378.06 ;
     RECT  635.14 515.24 641.86 515.44 ;
     RECT  641.86 365.68 642.62 378.06 ;
     RECT  638.78 260.26 642.82 264.66 ;
     RECT  635.62 176.68 643.3 176.88 ;
     RECT  635.14 529.1 643.3 529.3 ;
     RECT  632.74 275.38 643.78 285.24 ;
     RECT  642.62 365.68 644.74 381.42 ;
     RECT  630.34 566.06 645.02 566.26 ;
     RECT  645.02 566.06 645.7 572.98 ;
     RECT  645.7 572.78 646.18 572.98 ;
     RECT  644.74 373.66 647.14 381.42 ;
     RECT  624.58 666.86 647.14 693.52 ;
     RECT  642.82 264.04 647.62 264.66 ;
     RECT  641.86 349.72 647.9 355.38 ;
     RECT  641.86 331.66 648.58 335.64 ;
     RECT  647.14 373.66 648.58 373.86 ;
     RECT  647.14 673.16 648.58 693.52 ;
     RECT  647.9 347.2 650.5 355.38 ;
     RECT  650.5 347.2 650.98 354.96 ;
     RECT  648.58 673.16 650.98 687.64 ;
     RECT  643.78 275.38 651.46 275.58 ;
     RECT  650.98 347.2 652.9 347.4 ;
     RECT  638.5 644.18 653.38 644.38 ;
     RECT  646.94 290.08 654.34 294.48 ;
     RECT  641.66 312.76 654.34 317.16 ;
     RECT  647.62 264.46 655.3 264.66 ;
     RECT  648.58 331.66 655.3 332.28 ;
     RECT  652.7 233.38 655.78 233.58 ;
     RECT  655.3 332.08 656.26 332.28 ;
     RECT  648.86 158.2 657.22 158.4 ;
     RECT  650.98 680.3 658.18 687.64 ;
     RECT  654.34 316.96 660.58 317.16 ;
     RECT  654.34 290.08 661.06 290.28 ;
     RECT  658.18 687.44 668.74 687.64 ;
     RECT  655.58 595.04 670.18 595.24 ;
    LAYER Metal5 ;
     RECT  182.3 137.24 182.5 137.66 ;
     RECT  255.26 130.52 255.46 138.08 ;
     RECT  241.82 137.24 242.02 138.92 ;
     RECT  255.26 138.08 256.42 138.92 ;
     RECT  241.82 138.92 256.42 145.64 ;
     RECT  240.38 145.64 256.42 149 ;
     RECT  165.02 142.7 165.22 150.26 ;
     RECT  165.02 150.26 170.98 152.36 ;
     RECT  182.3 137.66 186.82 152.36 ;
     RECT  152.06 157.82 152.26 159.92 ;
     RECT  209.18 156.56 209.38 163.28 ;
     RECT  231.26 149 256.42 164.54 ;
     RECT  223.58 164.54 256.42 165.8 ;
     RECT  145.34 159.92 152.26 167.48 ;
     RECT  221.66 165.8 256.42 171.26 ;
     RECT  202.94 163.28 209.38 172.1 ;
     RECT  219.74 171.26 256.42 172.1 ;
     RECT  165.02 152.36 186.82 189.74 ;
     RECT  145.34 167.48 152.74 191.42 ;
     RECT  138.14 191.42 152.74 195.62 ;
     RECT  202.94 172.1 256.42 199.4 ;
     RECT  270.14 147.32 270.34 199.4 ;
     RECT  202.94 199.4 270.34 201.7 ;
     RECT  135.74 195.62 152.74 218.3 ;
     RECT  165.02 189.74 190.66 221.24 ;
     RECT  202.94 201.7 208.42 239.72 ;
     RECT  218.78 201.7 270.34 239.72 ;
     RECT  97.82 149.42 98.02 243.5 ;
     RECT  165.02 221.24 192.1 251.48 ;
     RECT  202.94 239.72 270.34 251.48 ;
     RECT  121.82 246.86 122.02 251.9 ;
     RECT  135.26 218.3 152.74 251.9 ;
     RECT  88.7 243.5 98.02 274.16 ;
     RECT  121.82 251.9 152.74 277.52 ;
     RECT  77.18 244.34 77.38 277.94 ;
     RECT  88.7 274.16 105.7 277.94 ;
     RECT  121.82 277.52 153.7 279.2 ;
     RECT  77.18 277.94 105.7 281.92 ;
     RECT  121.82 279.2 155.14 285.08 ;
     RECT  165.02 251.48 270.34 292.22 ;
     RECT  79.1 281.92 105.7 302.3 ;
     RECT  116.54 285.08 155.14 302.3 ;
     RECT  79.1 302.3 155.14 309.02 ;
     RECT  73.34 309.02 155.14 330.64 ;
     RECT  116.54 330.64 155.14 343.04 ;
     RECT  165.02 292.22 276.1 343.04 ;
     RECT  33.98 292.22 34.18 356.26 ;
     RECT  73.34 330.64 105.7 360.68 ;
     RECT  313.82 359 314.02 363.62 ;
     RECT  116.54 343.04 276.1 363.82 ;
     RECT  313.82 363.62 314.98 364.04 ;
     RECT  313.82 364.04 316.42 368.66 ;
     RECT  117.02 363.82 276.1 372.22 ;
     RECT  49.34 280.88 49.54 377.48 ;
     RECT  130.94 372.22 276.1 381.68 ;
     RECT  130.94 381.68 284.26 382.1 ;
     RECT  117.02 372.22 120.58 383.36 ;
     RECT  130.94 382.1 285.22 383.36 ;
     RECT  313.34 368.66 316.42 385.04 ;
     RECT  303.74 385.04 316.42 385.88 ;
     RECT  36.86 364.88 37.06 387.76 ;
     RECT  298.46 385.88 316.42 388.82 ;
     RECT  117.02 383.36 285.22 391.76 ;
     RECT  297.98 388.82 316.42 391.76 ;
     RECT  48.86 377.48 49.54 392.18 ;
     RECT  346.46 392.6 346.66 393.02 ;
     RECT  117.02 391.76 316.42 393.44 ;
     RECT  327.26 366.14 327.46 393.44 ;
     RECT  39.74 392.18 49.54 402.88 ;
     RECT  346.46 393.02 349.06 403.52 ;
     RECT  370.46 401 370.66 406.88 ;
     RECT  385.34 406.46 385.54 406.88 ;
     RECT  44.54 402.88 49.54 413.18 ;
     RECT  65.18 360.68 105.7 413.18 ;
     RECT  346.46 403.52 356.26 414.02 ;
     RECT  370.46 406.88 385.54 414.02 ;
     RECT  346.46 414.02 385.54 414.44 ;
     RECT  44.54 413.18 105.7 421.16 ;
     RECT  117.02 393.44 327.46 421.16 ;
     RECT  346.46 414.44 392.74 434.18 ;
     RECT  422.3 431.66 422.5 434.6 ;
     RECT  538.94 433.76 539.14 434.6 ;
     RECT  484.7 431.66 484.9 435.02 ;
     RECT  346.46 434.18 396.1 435.44 ;
     RECT  538.94 434.6 540.58 435.44 ;
     RECT  420.86 434.6 422.5 435.86 ;
     RECT  484.7 435.02 490.18 435.86 ;
     RECT  413.66 435.86 425.38 436.28 ;
     RECT  437.18 433.76 437.38 436.28 ;
     RECT  504.38 434.18 504.58 436.28 ;
     RECT  484.7 435.86 490.66 436.7 ;
     RECT  504.38 436.28 513.22 436.7 ;
     RECT  346.46 435.44 398.98 437.12 ;
     RECT  413.66 436.28 437.38 437.54 ;
     RECT  484.7 436.7 513.22 437.54 ;
     RECT  346.46 437.12 401.86 440.06 ;
     RECT  413.66 437.54 446.5 440.06 ;
     RECT  538.94 435.44 546.34 441.1 ;
     RECT  468.38 440.06 468.58 441.4 ;
     RECT  346.46 440.06 446.5 441.94 ;
     RECT  467.42 441.4 468.58 442.16 ;
     RECT  484.7 437.54 519.46 442.36 ;
     RECT  484.7 442.36 493.54 443.62 ;
     RECT  467.42 442.16 469.54 443.68 ;
     RECT  346.46 441.94 401.86 444.04 ;
     RECT  484.7 443.62 492.1 444.26 ;
     RECT  464.06 443.68 469.54 446.14 ;
     RECT  346.46 444.04 398.98 446.98 ;
     RECT  464.06 446.14 469.06 447.2 ;
     RECT  481.34 444.26 492.1 447.2 ;
     RECT  413.66 441.94 446.5 448.24 ;
     RECT  431.42 448.24 446.5 448.46 ;
     RECT  460.22 447.2 469.06 448.46 ;
     RECT  510.62 442.36 519.46 449.72 ;
     RECT  431.42 448.46 469.06 450.34 ;
     RECT  44.54 421.16 327.46 451.6 ;
     RECT  546.62 451.82 546.82 452.24 ;
     RECT  510.62 449.72 523.78 452.44 ;
     RECT  448.7 450.34 469.06 453.28 ;
     RECT  480.38 447.2 492.1 454.76 ;
     RECT  44.54 451.6 86.98 455.38 ;
     RECT  543.74 452.24 546.82 456.22 ;
     RECT  480.38 454.76 494.98 456.44 ;
     RECT  543.74 456.22 543.94 458.32 ;
     RECT  448.7 453.28 466.66 460.64 ;
     RECT  477.5 456.44 494.98 461.26 ;
     RECT  431.42 450.34 431.62 461.48 ;
     RECT  348.86 446.98 398.98 462.32 ;
     RECT  413.66 448.24 413.86 462.32 ;
     RECT  429.5 461.48 431.62 462.74 ;
     RECT  444.38 460.64 466.66 462.74 ;
     RECT  515.42 452.44 517.06 466.1 ;
     RECT  348.86 462.32 413.86 466.52 ;
     RECT  571.1 461.9 571.3 466.52 ;
     RECT  582.62 463.58 582.82 466.52 ;
     RECT  429.5 462.74 466.66 469.88 ;
     RECT  429.5 469.88 468.58 470.3 ;
     RECT  505.34 462.74 505.54 471.56 ;
     RECT  515.42 466.1 522.34 471.56 ;
     RECT  560.06 466.94 560.26 471.56 ;
     RECT  571.1 466.52 582.82 471.56 ;
     RECT  426.14 470.3 468.58 472.4 ;
     RECT  480.38 461.26 494.98 474.08 ;
     RECT  96.86 451.6 327.46 474.92 ;
     RECT  340.22 466.52 413.86 474.92 ;
     RECT  479.9 474.08 494.98 474.92 ;
     RECT  505.34 471.56 522.34 474.92 ;
     RECT  560.06 471.56 582.82 474.92 ;
     RECT  45.5 455.38 86.98 477.22 ;
     RECT  552.86 474.92 582.82 477.44 ;
     RECT  545.66 477.44 582.82 478.06 ;
     RECT  96.86 474.92 413.86 480.8 ;
     RECT  426.14 472.4 469.06 480.8 ;
     RECT  545.66 478.06 576.58 482.06 ;
     RECT  538.94 482.06 576.58 485.62 ;
     RECT  96.86 480.8 469.06 485.84 ;
     RECT  479.9 474.92 522.34 485.84 ;
     RECT  550.94 485.62 571.3 488.56 ;
     RECT  538.94 485.62 540.1 494.02 ;
     RECT  45.5 477.22 75.46 496.54 ;
     RECT  550.94 488.56 566.02 500.74 ;
     RECT  86.78 477.22 86.98 504.1 ;
     RECT  550.94 500.74 562.18 508.72 ;
     RECT  96.86 485.84 522.34 508.94 ;
     RECT  96.86 508.94 527.14 529.52 ;
     RECT  538.94 494.02 539.14 531.2 ;
     RECT  550.94 508.72 557.86 531.2 ;
     RECT  538.94 531.2 557.86 533.72 ;
     RECT  45.5 496.54 72.1 538.54 ;
     RECT  47.9 538.54 72.1 539.8 ;
     RECT  96.86 529.52 529.06 545.48 ;
     RECT  538.94 533.72 565.06 545.48 ;
     RECT  96.86 545.48 569.86 554.3 ;
     RECT  55.58 539.8 72.1 556.6 ;
     RECT  58.46 556.6 72.1 557.44 ;
     RECT  96.86 554.3 578.98 559.34 ;
     RECT  590.78 555.14 590.98 559.34 ;
     RECT  29.66 409.4 29.86 561.64 ;
     RECT  96.86 559.34 590.98 562.48 ;
     RECT  143.42 562.48 590.98 564.8 ;
     RECT  67.1 557.44 72.1 576.76 ;
     RECT  143.42 564.8 592.9 576.76 ;
     RECT  67.1 576.76 71.14 579.28 ;
     RECT  143.42 576.76 590.98 582.22 ;
     RECT  143.42 582.22 583.3 583.9 ;
     RECT  143.42 583.9 327.94 586 ;
     RECT  144.86 586 327.94 587.68 ;
     RECT  67.1 579.28 67.3 591.88 ;
     RECT  209.66 587.68 327.94 598.4 ;
     RECT  341.18 583.9 583.3 598.6 ;
     RECT  144.86 587.68 197.86 599.44 ;
     RECT  96.86 562.48 133.54 601.96 ;
     RECT  144.86 599.44 180.58 602.8 ;
     RECT  209.66 598.4 329.38 604.9 ;
     RECT  341.18 598.6 575.62 604.9 ;
     RECT  341.18 604.9 534.82 605.74 ;
     RECT  553.82 604.9 575.62 605.74 ;
     RECT  553.82 605.74 557.86 606.16 ;
     RECT  571.1 605.74 575.62 606.58 ;
     RECT  534.62 605.74 534.82 607 ;
     RECT  216.38 604.9 329.38 608.06 ;
     RECT  341.18 605.74 521.38 608.06 ;
     RECT  105.02 601.96 133.54 609.52 ;
     RECT  575.42 606.58 575.62 610.36 ;
     RECT  216.38 608.06 521.38 611.62 ;
     RECT  553.82 606.16 554.02 612.88 ;
     RECT  105.02 609.52 127.3 613.3 ;
     RECT  341.18 611.62 521.38 613.3 ;
     RECT  154.46 602.8 180.58 614.98 ;
     RECT  105.02 613.3 122.02 617.92 ;
     RECT  115.58 617.92 122.02 618.34 ;
     RECT  341.18 613.3 454.18 621.92 ;
     RECT  216.38 611.62 329.38 625.48 ;
     RECT  216.38 625.48 216.58 632.2 ;
     RECT  339.74 621.92 454.18 632.62 ;
     RECT  230.78 625.48 329.38 633.04 ;
     RECT  339.74 632.62 339.94 633.46 ;
     RECT  119.9 618.34 122.02 647.74 ;
     RECT  119.9 647.74 120.1 651.1 ;
     RECT  190.46 599.44 197.86 652.36 ;
     RECT  105.02 617.92 105.22 654.88 ;
     RECT  352.7 632.62 454.18 655.72 ;
     RECT  154.46 614.98 176.26 673.36 ;
     RECT  468.38 613.3 521.38 673.78 ;
     RECT  230.78 633.04 277.06 680.5 ;
     RECT  270.14 680.5 277.06 688.48 ;
     RECT  230.78 680.5 255.94 688.9 ;
     RECT  190.46 652.36 193.06 689.32 ;
     RECT  468.38 673.78 473.38 689.74 ;
     RECT  353.18 655.72 454.18 691.42 ;
     RECT  471.74 689.74 473.38 691.42 ;
     RECT  485.66 673.78 521.38 691.42 ;
     RECT  471.74 691.42 471.94 692.68 ;
     RECT  514.94 691.42 521.38 693.1 ;
     RECT  230.78 688.9 250.18 693.52 ;
     RECT  271.58 688.48 277.06 693.52 ;
     RECT  385.34 691.42 392.74 693.94 ;
     RECT  515.9 693.1 521.38 693.94 ;
     RECT  413.66 691.42 422.98 694.36 ;
     RECT  154.46 673.36 154.66 694.78 ;
     RECT  413.66 694.36 413.86 694.78 ;
     RECT  230.78 693.52 235.78 695.2 ;
     RECT  291.74 633.04 329.38 695.2 ;
     RECT  353.18 691.42 373.54 695.2 ;
     RECT  521.18 693.94 521.38 695.2 ;
     RECT  370.46 695.2 373.54 695.62 ;
     RECT  191.42 689.32 193.06 696.04 ;
     RECT  370.46 695.62 371.62 696.04 ;
     RECT  169.34 673.36 176.26 696.46 ;
     RECT  370.46 696.04 370.66 696.46 ;
     RECT  169.34 696.46 171.46 696.88 ;
     RECT  291.74 695.2 306.82 696.88 ;
     RECT  385.34 693.94 385.54 696.88 ;
     RECT  169.34 696.88 170.5 697.3 ;
     RECT  298.46 696.88 306.82 697.3 ;
     RECT  169.34 697.3 169.54 697.72 ;
     RECT  298.46 697.3 298.66 697.72 ;
     RECT  485.66 691.42 485.86 698.14 ;
     RECT  248.06 693.52 248.26 698.56 ;
     RECT  191.42 696.04 191.62 698.98 ;
  END
END core_wrap
END LIBRARY
