VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA croc_chip_via1_2_10000_440_1_24_410_410
  VIARULE via1Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.01 0.125 0.05 0.005 ;
  ROWCOL 1 24 ;
END croc_chip_via1_2_10000_440_1_24_410_410

VIA croc_chip_via2_3_10000_200_1_24_410_410
  VIARULE via2Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 24 ;
END croc_chip_via2_3_10000_200_1_24_410_410

VIA croc_chip_via3_4_10000_200_1_24_410_410
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.005 0.05 0.05 0.005 ;
  ROWCOL 1 24 ;
END croc_chip_via3_4_10000_200_1_24_410_410

VIA croc_chip_via4_5_10000_200_1_24_410_410
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 24 ;
END croc_chip_via4_5_10000_200_1_24_410_410

VIA croc_chip_via5_6_10000_1500_1_11_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.42 ;
  ROWCOL 1 11 ;
END croc_chip_via5_6_10000_1500_1_11_840_840

VIA croc_chip_via6_7_10000_2860_1_5_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.5 0.63 0.5 ;
  ROWCOL 1 5 ;
END croc_chip_via6_7_10000_2860_1_5_1960_1960

VIA croc_chip_via1_2_6000_440_1_14_410_410
  VIARULE via1Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.01 0.125 0.05 0.005 ;
  ROWCOL 1 14 ;
END croc_chip_via1_2_6000_440_1_14_410_410

VIA croc_chip_via2_3_6000_200_1_14_410_410
  VIARULE via2Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 14 ;
END croc_chip_via2_3_6000_200_1_14_410_410

VIA croc_chip_via3_4_6000_200_1_14_410_410
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.005 0.05 0.05 0.005 ;
  ROWCOL 1 14 ;
END croc_chip_via3_4_6000_200_1_14_410_410

VIA croc_chip_via4_5_6000_200_1_14_410_410
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 14 ;
END croc_chip_via4_5_6000_200_1_14_410_410

VIA croc_chip_via5_6_6000_1500_1_6_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.42 ;
  ROWCOL 1 6 ;
END croc_chip_via5_6_6000_1500_1_6_840_840

VIA croc_chip_via6_7_6000_2860_1_3_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.5 0.59 0.5 ;
  ROWCOL 1 3 ;
END croc_chip_via6_7_6000_2860_1_3_1960_1960

VIA croc_chip_via1_2_2000_440_1_5_410_410
  VIARULE via1Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.01 0.125 0.05 0.005 ;
  ROWCOL 1 5 ;
END croc_chip_via1_2_2000_440_1_5_410_410

VIA croc_chip_via2_3_2000_200_1_5_410_410
  VIARULE via2Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 5 ;
END croc_chip_via2_3_2000_200_1_5_410_410

VIA croc_chip_via3_4_2000_200_1_5_410_410
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.005 0.05 0.05 0.005 ;
  ROWCOL 1 5 ;
END croc_chip_via3_4_2000_200_1_5_410_410

VIA croc_chip_via4_5_2000_200_1_5_410_410
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 5 ;
END croc_chip_via4_5_2000_200_1_5_410_410

VIA croc_chip_via5_6_2000_1500_1_1_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.42 ;
END croc_chip_via5_6_2000_1500_1_1_840_840

VIA croc_chip_via6_7_2000_1650_1_1_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.5 0.55 0.5 ;
END croc_chip_via6_7_2000_1650_1_1_1960_1960

VIA croc_chip_via1_2_1880_440_1_4_410_410
  VIARULE via1Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.01 0.125 0.05 0.005 ;
  ROWCOL 1 4 ;
END croc_chip_via1_2_1880_440_1_4_410_410

VIA croc_chip_via2_3_1880_760_1_4_480_480
  VIARULE via2Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 4 ;
END croc_chip_via2_3_1880_760_1_4_480_480

VIA croc_chip_via3_4_1880_760_1_4_480_480
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.005 0.05 0.05 0.005 ;
  ROWCOL 1 4 ;
END croc_chip_via3_4_1880_760_1_4_480_480

VIA croc_chip_via4_5_1880_760_1_4_480_480
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 4 ;
END croc_chip_via4_5_1880_760_1_4_480_480

VIA croc_chip_via5_6_1880_1500_1_1_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.42 ;
END croc_chip_via5_6_1880_1500_1_1_840_840

VIA croc_chip_via6_7_10000_10000_5_5_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.63 0.5 ;
  ROWCOL 5 5 ;
END croc_chip_via6_7_10000_10000_5_5_1960_1960

VIA croc_chip_via6_7_13330_18000_9_6_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 1.315 0.71 1.315 0.5 ;
  ROWCOL 9 6 ;
END croc_chip_via6_7_13330_18000_9_6_1960_1960

VIA croc_chip_via6_7_13330_10000_5_6_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 1.315 0.5 ;
  ROWCOL 5 6 ;
END croc_chip_via6_7_13330_10000_5_6_1960_1960

VIA croc_chip_via6_7_20000_10000_5_10_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.73 0.5 ;
  ROWCOL 5 10 ;
END croc_chip_via6_7_20000_10000_5_10_1960_1960

VIA croc_chip_via6_7_20000_18000_9_10_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.73 0.71 0.73 0.5 ;
  ROWCOL 9 10 ;
END croc_chip_via6_7_20000_18000_9_10_1960_1960

VIA croc_chip_via6_7_6000_10000_5_3_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.59 0.5 ;
  ROWCOL 5 3 ;
END croc_chip_via6_7_6000_10000_5_3_1960_1960

VIA croc_chip_via2_3_2000_440_1_5_410_410
  VIARULE via2Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.085 0.05 ;
  ROWCOL 1 5 ;
END croc_chip_via2_3_2000_440_1_5_410_410

VIA croc_chip_via3_4_2000_2000_4_4_480_480
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.185 0.05 0.05 0.185 ;
  ROWCOL 4 4 ;
END croc_chip_via3_4_2000_2000_4_4_480_480

VIA croc_chip_via3_4_2000_6000_12_4_480_480
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.185 0.05 0.05 0.005 ;
  ROWCOL 12 4 ;
END croc_chip_via3_4_2000_6000_12_4_480_480

VIA croc_chip_via4_5_2000_6000_12_4_480_480
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 12 4 ;
END croc_chip_via4_5_2000_6000_12_4_480_480

VIA croc_chip_via5_6_2000_6000_6_1_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.69 ;
  ROWCOL 6 1 ;
END croc_chip_via5_6_2000_6000_6_1_840_840

VIA croc_chip_via4_5_2810_6000_12_6_480_480
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.11 0.265 0.005 0.05 ;
  ROWCOL 12 6 ;
END croc_chip_via4_5_2810_6000_12_6_480_480

VIA croc_chip_via5_6_2810_6000_6_2_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.69 ;
  ROWCOL 6 2 ;
END croc_chip_via5_6_2810_6000_6_2_840_840

VIA croc_chip_via6_7_6000_6000_3_3_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.59 0.59 0.5 ;
  ROWCOL 3 3 ;
END croc_chip_via6_7_6000_6000_3_3_1960_1960

MACRO croc_chip
  FOREIGN croc_chip 0 0 ;
  CLASS BLOCK ;
  SIZE 1870 BY 1870 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 997 0 1067 ;
    END
  END clk_i
  PIN fetch_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1173 0 1243 ;
    END
  END fetch_en_i
  PIN gpio0_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  381 -70 451 0 ;
    END
  END gpio0_io
  PIN gpio10_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1261 -70 1331 0 ;
    END
  END gpio10_io
  PIN gpio11_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1349 -70 1419 0 ;
    END
  END gpio11_io
  PIN gpio12_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 381 1870 451 ;
    END
  END gpio12_io
  PIN gpio13_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 469 1870 539 ;
    END
  END gpio13_io
  PIN gpio14_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 557 1870 627 ;
    END
  END gpio14_io
  PIN gpio15_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 645 1870 715 ;
    END
  END gpio15_io
  PIN gpio16_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 733 1870 803 ;
    END
  END gpio16_io
  PIN gpio17_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 821 1870 891 ;
    END
  END gpio17_io
  PIN gpio18_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 909 1870 979 ;
    END
  END gpio18_io
  PIN gpio19_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 997 1870 1067 ;
    END
  END gpio19_io
  PIN gpio1_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  469 -70 539 0 ;
    END
  END gpio1_io
  PIN gpio20_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 1085 1870 1155 ;
    END
  END gpio20_io
  PIN gpio21_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 1173 1870 1243 ;
    END
  END gpio21_io
  PIN gpio22_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 1261 1870 1331 ;
    END
  END gpio22_io
  PIN gpio23_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1800 1349 1870 1419 ;
    END
  END gpio23_io
  PIN gpio24_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1349 1800 1419 1870 ;
    END
  END gpio24_io
  PIN gpio25_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1261 1800 1331 1870 ;
    END
  END gpio25_io
  PIN gpio26_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1173 1800 1243 1870 ;
    END
  END gpio26_io
  PIN gpio27_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1085 1800 1155 1870 ;
    END
  END gpio27_io
  PIN gpio28_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  997 1800 1067 1870 ;
    END
  END gpio28_io
  PIN gpio29_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  909 1800 979 1870 ;
    END
  END gpio29_io
  PIN gpio2_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  557 -70 627 0 ;
    END
  END gpio2_io
  PIN gpio30_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  821 1800 891 1870 ;
    END
  END gpio30_io
  PIN gpio31_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  733 1800 803 1870 ;
    END
  END gpio31_io
  PIN gpio3_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  645 -70 715 0 ;
    END
  END gpio3_io
  PIN gpio4_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  733 -70 803 0 ;
    END
  END gpio4_io
  PIN gpio5_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  821 -70 891 0 ;
    END
  END gpio5_io
  PIN gpio6_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  909 -70 979 0 ;
    END
  END gpio6_io
  PIN gpio7_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  997 -70 1067 0 ;
    END
  END gpio7_io
  PIN gpio8_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1085 -70 1155 0 ;
    END
  END gpio8_io
  PIN gpio9_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1173 -70 1243 0 ;
    END
  END gpio9_io
  PIN jtag_tck_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 733 0 803 ;
    END
  END jtag_tck_i
  PIN jtag_tdi_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 469 0 539 ;
    END
  END jtag_tdi_i
  PIN jtag_tdo_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 381 0 451 ;
    END
  END jtag_tdo_o
  PIN jtag_tms_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 557 0 627 ;
    END
  END jtag_tms_i
  PIN jtag_trst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 645 0 715 ;
    END
  END jtag_trst_ni
  PIN ref_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 909 0 979 ;
    END
  END ref_clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 821 0 891 ;
    END
  END rst_ni
  PIN status_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1085 0 1155 ;
    END
  END status_o
  PIN uart_rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1349 0 1419 ;
    END
  END uart_rx_i
  PIN uart_tx_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1261 0 1331 ;
    END
  END uart_tx_o
  PIN unused0_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  645 1800 715 1870 ;
    END
  END unused0_o
  PIN unused1_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  557 1800 627 1870 ;
    END
  END unused1_o
  PIN unused2_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  469 1800 539 1870 ;
    END
  END unused2_o
  PIN unused3_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  381 1800 451 1870 ;
    END
  END unused3_o
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER TopMetal2 ;
        RECT  205 1800 275 1870 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  1800 1525 1870 1595 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  1525 -70 1595 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 205 0 275 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER TopMetal2 ;
        RECT  1437 1800 1507 1870 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  1800 293 1870 363 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  293 -70 363 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1437 0 1507 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal2 ;
        RECT  293 1800 363 1870 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  1800 1437 1870 1507 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  1437 -70 1507 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 293 0 363 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal2 ;
        RECT  1525 1800 1595 1870 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  1800 205 1870 275 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  205 -70 275 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1525 0 1595 ;
    END
  END VSSIO
  OBS
    LAYER Metal1 ;
     RECT  205 -70 275 0 ;
     RECT  293 -70 363 0 ;
     RECT  381 -70 451 0 ;
     RECT  469 -70 539 0 ;
     RECT  557 -70 627 0 ;
     RECT  645 -70 715 0 ;
     RECT  733 -70 803 0 ;
     RECT  821 -70 891 0 ;
     RECT  909 -70 979 0 ;
     RECT  997 -70 1067 0 ;
     RECT  1085 -70 1155 0 ;
     RECT  1173 -70 1243 0 ;
     RECT  1261 -70 1331 0 ;
     RECT  1349 -70 1419 0 ;
     RECT  1437 -70 1507 0 ;
     RECT  1525 -70 1595 0 ;
     RECT  0 0 1800 180 ;
     RECT  0 180 180 205 ;
     RECT  1620 180 1800 205 ;
     RECT  -70 205 180 219.02 ;
     RECT  202 215.24 1598 219.02 ;
     RECT  1620 205 1870 219.02 ;
     RECT  -70 219.02 1870 275 ;
     RECT  0 275 1800 293 ;
     RECT  -70 293 1870 363 ;
     RECT  0 363 1800 381 ;
     RECT  -70 381 1870 451 ;
     RECT  0 451 1800 469 ;
     RECT  -70 469 1870 539 ;
     RECT  0 539 1800 557 ;
     RECT  -70 557 1870 627 ;
     RECT  0 627 1800 645 ;
     RECT  -70 645 1870 715 ;
     RECT  0 715 1800 733 ;
     RECT  -70 733 1870 803 ;
     RECT  0 803 1800 821 ;
     RECT  -70 821 1870 877.18 ;
     RECT  -70 877.18 217.44 891 ;
     RECT  897.12 877.18 1870 891 ;
     RECT  897.12 891 1800 905.76 ;
     RECT  0 891 217.44 909 ;
     RECT  245.28 905.76 1800 909 ;
     RECT  -70 909 217.44 979 ;
     RECT  245.28 909 1870 979 ;
     RECT  0 979 217.44 997 ;
     RECT  245.28 979 1800 997 ;
     RECT  -70 997 217.44 1067 ;
     RECT  245.28 997 1870 1067 ;
     RECT  0 1067 217.44 1085 ;
     RECT  245.28 1067 1800 1085 ;
     RECT  -70 1085 217.44 1155 ;
     RECT  245.28 1085 1870 1155 ;
     RECT  0 1155 217.44 1173 ;
     RECT  245.28 1155 1800 1173 ;
     RECT  -70 1173 217.44 1243 ;
     RECT  245.28 1173 1870 1243 ;
     RECT  0 1243 217.44 1261 ;
     RECT  245.28 1243 1800 1261 ;
     RECT  -70 1261 217.44 1331 ;
     RECT  245.28 1261 1870 1331 ;
     RECT  0 1331 217.44 1349 ;
     RECT  245.28 1331 1800 1349 ;
     RECT  245.28 1349 1870 1372.36 ;
     RECT  245.28 1372.36 903.84 1382 ;
     RECT  1114.08 1372.36 1870 1382 ;
     RECT  -70 1349 217.44 1419 ;
     RECT  245.28 1382 1870 1419 ;
     RECT  0 1419 217.44 1437 ;
     RECT  245.28 1419 1800 1437 ;
     RECT  -70 1437 217.44 1507 ;
     RECT  245.28 1437 1870 1507 ;
     RECT  0 1507 217.44 1525 ;
     RECT  245.28 1507 1800 1525 ;
     RECT  245.28 1525 1870 1552.58 ;
     RECT  -70 1525 217.44 1579.82 ;
     RECT  897.12 1552.58 1870 1579.82 ;
     RECT  -70 1579.82 1870 1580.26 ;
     RECT  202 1580.26 1598 1584.04 ;
     RECT  -70 1580.26 180 1595 ;
     RECT  1620 1580.26 1870 1595 ;
     RECT  0 1595 180 1620 ;
     RECT  1620 1595 1800 1620 ;
     RECT  0 1620 1800 1800 ;
     RECT  205 1800 275 1870 ;
     RECT  293 1800 363 1870 ;
     RECT  381 1800 451 1870 ;
     RECT  469 1800 539 1870 ;
     RECT  557 1800 627 1870 ;
     RECT  645 1800 715 1870 ;
     RECT  733 1800 803 1870 ;
     RECT  821 1800 891 1870 ;
     RECT  909 1800 979 1870 ;
     RECT  997 1800 1067 1870 ;
     RECT  1085 1800 1155 1870 ;
     RECT  1173 1800 1243 1870 ;
     RECT  1261 1800 1331 1870 ;
     RECT  1349 1800 1419 1870 ;
     RECT  1437 1800 1507 1870 ;
     RECT  1525 1800 1595 1870 ;
    LAYER Metal2 ;
     RECT  -70 205 0 275 ;
     RECT  -70 293 0 363 ;
     RECT  -70 381 0 451 ;
     RECT  -70 469 0 539 ;
     RECT  -70 557 0 627 ;
     RECT  -70 645 0 715 ;
     RECT  -70 733 0 803 ;
     RECT  -70 821 0 891 ;
     RECT  -70 909 0 979 ;
     RECT  -70 997 0 1067 ;
     RECT  -70 1085 0 1155 ;
     RECT  -70 1173 0 1243 ;
     RECT  -70 1261 0 1331 ;
     RECT  -70 1349 0 1419 ;
     RECT  -70 1437 0 1507 ;
     RECT  -70 1525 0 1595 ;
     RECT  0 0 180 1800 ;
     RECT  180 219.14 202.14 1580.14 ;
     RECT  180 0 205 180 ;
     RECT  180 1620 205 1800 ;
     RECT  202.14 215.36 211.86 1583.92 ;
     RECT  211.86 423.26 215.005 549.04 ;
     RECT  211.86 701.3 215.005 831.7 ;
     RECT  211.86 1117.94 216.1 1118.98 ;
     RECT  215.005 427.04 217.605 549.04 ;
     RECT  216.1 1118.78 219.46 1118.98 ;
     RECT  211.86 874.75 223.235 875.815 ;
     RECT  217.605 427.35 223.34 549.04 ;
     RECT  223.235 874.75 223.685 874.98 ;
     RECT  223.34 427.35 229.34 549.88 ;
     RECT  229.34 424.1 229.82 549.88 ;
     RECT  229.82 420.32 230.02 549.88 ;
     RECT  227.42 1565.66 233.66 1565.86 ;
     RECT  215.005 701.3 234.62 828.03 ;
     RECT  230.02 423.26 235.1 549.88 ;
     RECT  235.1 423.26 235.58 553.66 ;
     RECT  223.685 874.76 236.06 874.96 ;
     RECT  236.06 874.76 236.54 875.8 ;
     RECT  229.82 1577.42 237.5 1577.62 ;
     RECT  237.5 1577.42 239.42 1578.04 ;
     RECT  240.86 837.38 241.34 837.58 ;
     RECT  235.58 423.26 241.82 554.92 ;
     RECT  236.54 874.76 242.3 877.48 ;
     RECT  234.62 697.52 242.78 828.03 ;
     RECT  241.34 836.54 242.78 837.58 ;
     RECT  242.78 697.52 243.26 837.58 ;
     RECT  242.3 869.3 243.26 877.48 ;
     RECT  241.82 423.26 243.74 555.34 ;
     RECT  243.26 869.3 243.74 877.9 ;
     RECT  243.74 423.26 245.18 556.6 ;
     RECT  243.26 693.74 245.18 837.58 ;
     RECT  245.18 1218.36 245.575 1221.5 ;
     RECT  245.18 1240.62 245.575 1240.82 ;
     RECT  245.575 1032.3 245.66 1032.5 ;
     RECT  245.575 1130.16 245.66 1130.36 ;
     RECT  245.575 1210.38 245.66 1221.5 ;
     RECT  245.575 1233.06 245.66 1240.82 ;
     RECT  245.575 1263.72 245.66 1271.48 ;
     RECT  245.575 1301.1 245.66 1309.28 ;
     RECT  245.575 999.12 246.055 1006.88 ;
     RECT  245.575 1021.8 246.055 1022 ;
     RECT  245.66 1263.72 246.055 1281.14 ;
     RECT  245.66 1123.02 246.14 1130.36 ;
     RECT  245.575 1160.4 246.14 1160.6 ;
     RECT  245.575 1173 246.14 1173.2 ;
     RECT  245.66 1202.82 246.14 1221.5 ;
     RECT  245.66 1230.12 246.14 1240.82 ;
     RECT  246.055 1258.68 246.14 1281.14 ;
     RECT  246.055 999.12 246.355 1022 ;
     RECT  245.575 1062.12 246.355 1069.88 ;
     RECT  246.14 1122.6 246.355 1130.36 ;
     RECT  245.575 1145.28 246.355 1145.48 ;
     RECT  245.575 1188.12 246.355 1188.32 ;
     RECT  245.575 1319.16 246.355 1319.36 ;
     RECT  245.575 1099.92 246.495 1105.16 ;
     RECT  245.66 1032.3 246.535 1033.34 ;
     RECT  246.14 1258.68 246.535 1289.12 ;
     RECT  245.66 1300.26 246.535 1309.28 ;
     RECT  246.14 1160.4 246.62 1173.2 ;
     RECT  246.535 1032.3 247.015 1039.64 ;
     RECT  246.355 1062.12 247.015 1070.72 ;
     RECT  246.62 1079.76 247.015 1082.06 ;
     RECT  246.14 1199.04 247.045 1242.08 ;
     RECT  247.015 1032.3 247.1 1044.68 ;
     RECT  246.62 1160.4 247.1 1176.14 ;
     RECT  247.045 1199.04 247.1 1248.8 ;
     RECT  246.535 1258.68 247.1 1309.28 ;
     RECT  246.355 1187.28 247.525 1188.32 ;
     RECT  247.1 1199.04 247.525 1309.28 ;
     RECT  247.1 1032.3 247.58 1052.66 ;
     RECT  247.015 1062.12 247.58 1082.06 ;
     RECT  246.495 1092.99 247.58 1105.16 ;
     RECT  247.58 1092.78 247.935 1105.16 ;
     RECT  247.58 1032.3 247.975 1082.06 ;
     RECT  247.935 1092.78 247.975 1112.09 ;
     RECT  246.355 1145.28 248.06 1146.32 ;
     RECT  246.355 1319.16 248.06 1320.2 ;
     RECT  245.18 420.32 248.54 556.6 ;
     RECT  247.975 1032.3 248.54 1112.09 ;
     RECT  246.355 1122.6 248.54 1131.2 ;
     RECT  248.06 1142.34 248.54 1146.32 ;
     RECT  247.1 1157.46 248.54 1177.82 ;
     RECT  247.525 1187.28 248.54 1309.28 ;
     RECT  248.06 1319.16 248.54 1321.46 ;
     RECT  248.54 1187.28 248.935 1322.72 ;
     RECT  246.355 998.28 249.02 1022 ;
     RECT  248.54 1031.04 249.02 1112.09 ;
     RECT  248.54 1122.6 249.415 1146.32 ;
     RECT  248.54 1157.46 249.415 1178.24 ;
     RECT  249.02 1031.04 249.5 1112.3 ;
     RECT  249.415 1122.6 249.5 1178.24 ;
     RECT  248.935 1187.28 249.715 1326.92 ;
     RECT  249.02 994.5 249.98 1022 ;
     RECT  249.5 1031.04 249.98 1178.24 ;
     RECT  249.715 1187.28 249.98 1327.76 ;
     RECT  245.18 693.32 250.46 837.58 ;
     RECT  250.46 1467.84 251.36 1468.04 ;
     RECT  249.98 994.5 252.295 1327.76 ;
     RECT  250.46 689.12 252.86 837.58 ;
     RECT  251.36 1466.83 252.86 1468.04 ;
     RECT  252.295 991.56 253.075 1327.76 ;
     RECT  252.86 1460.28 253.76 1468.04 ;
     RECT  254.3 1447.68 255.2 1447.88 ;
     RECT  248.54 416.96 255.74 556.6 ;
     RECT  255.2 1447.68 255.74 1448.89 ;
     RECT  253.76 1459.27 255.74 1468.04 ;
     RECT  252.86 687.44 257.18 837.58 ;
     RECT  255.74 410.24 258.62 556.6 ;
     RECT  258.62 410.24 259.3 557.86 ;
     RECT  259.015 978.96 259.795 979.16 ;
     RECT  259.795 978.96 259.975 980 ;
     RECT  253.075 990.72 260.06 1327.76 ;
     RECT  255.74 1447.68 260.06 1468.04 ;
     RECT  211.86 1479.56 260.06 1479.76 ;
     RECT  259.975 971.4 261.02 980 ;
     RECT  260.06 990.3 261.02 1327.76 ;
     RECT  261.02 971.4 262.22 1327.76 ;
     RECT  262.22 971.4 262.94 1331.12 ;
     RECT  259.3 410.24 263.9 556.18 ;
     RECT  260.06 1447.68 263.9 1479.76 ;
     RECT  243.74 869.3 264.32 878.32 ;
     RECT  262.94 971.4 264.38 1331.96 ;
     RECT  264.32 867.585 265.34 878.32 ;
     RECT  263.9 1447.26 265.82 1479.76 ;
     RECT  264.38 971.4 266.3 1334.48 ;
     RECT  265.82 1445.16 266.72 1479.76 ;
     RECT  266.3 971.4 267.26 1339.1 ;
     RECT  267.26 971.4 269.18 1342.46 ;
     RECT  235.58 857.54 270.08 857.74 ;
     RECT  265.34 867.2 270.08 878.32 ;
     RECT  269.18 971.4 270.62 1342.88 ;
     RECT  270.62 971.4 271.58 1343.3 ;
     RECT  266.72 1444.15 272.54 1479.76 ;
     RECT  211.86 388.4 273.5 388.6 ;
     RECT  271.58 968.46 273.98 1343.3 ;
     RECT  263.9 409.82 274.46 556.18 ;
     RECT  273.5 388.4 274.94 395.74 ;
     RECT  274.46 409.4 274.94 556.18 ;
     RECT  205 -70 275 180 ;
     RECT  205 1620 275 1870 ;
     RECT  273.98 966.78 277.255 1343.3 ;
     RECT  270.08 857.54 278.3 878.32 ;
     RECT  277.255 964.26 278.78 1343.3 ;
     RECT  255.26 615.62 279.74 615.82 ;
     RECT  279.625 1368.285 280.12 1368.515 ;
     RECT  272.54 1439.7 280.22 1479.76 ;
     RECT  278.3 856.28 280.9 878.32 ;
     RECT  280.22 1437.6 281.12 1479.76 ;
     RECT  281.12 1436.59 282.62 1479.76 ;
     RECT  282.62 1422.48 283.52 1479.76 ;
     RECT  278.78 964.26 283.61 1346.66 ;
     RECT  283.61 963.92 283.68 1346.66 ;
     RECT  283.58 1409.88 284.48 1410.08 ;
     RECT  274.94 388.4 285.5 556.18 ;
     RECT  284.48 1409.88 285.5 1411.09 ;
     RECT  283.52 1421.47 285.5 1479.76 ;
     RECT  283.68 963.84 286.49 1346.66 ;
     RECT  286.49 963.84 286.56 1347 ;
     RECT  285.5 388.4 286.94 557.02 ;
     RECT  286.56 963.84 289.34 1347.08 ;
     RECT  280.12 1368.285 289.82 1369.35 ;
     RECT  289.34 960.9 291.74 1347.08 ;
     RECT  275 0 293 180 ;
     RECT  275 1620 293 1800 ;
     RECT  289.82 1368.285 293.18 1369.76 ;
     RECT  285.5 1409.88 293.18 1479.76 ;
     RECT  293.18 1409.46 297.22 1479.76 ;
     RECT  291.74 956.28 298.94 1347.08 ;
     RECT  298.94 952.92 300.86 1347.08 ;
     RECT  300.86 946.2 301.76 1347.08 ;
     RECT  305.18 929.4 306.08 930.44 ;
     RECT  301.76 945.19 306.14 1347.08 ;
     RECT  293.18 1367.46 306.82 1369.76 ;
     RECT  306.08 929.4 307.1 930.475 ;
     RECT  297.22 1413.91 307.765 1479.76 ;
     RECT  306.14 942.84 308.425 1347.08 ;
     RECT  307.765 1415.34 310.18 1479.76 ;
     RECT  307.1 929.4 310.46 930.86 ;
     RECT  308.425 942.84 310.46 1350.875 ;
     RECT  310.18 1415.34 311.14 1430.66 ;
     RECT  286.94 388.4 311.19 557.86 ;
     RECT  279.74 615.62 311.19 616.66 ;
     RECT  211.86 629.9 311.19 630.1 ;
     RECT  301.82 651.32 311.19 651.52 ;
     RECT  293.66 673.16 311.19 673.36 ;
     RECT  257.18 684.5 311.19 837.58 ;
     RECT  280.9 857.54 311.19 878.32 ;
     RECT  239.42 1577 311.19 1578.04 ;
     RECT  310.46 926.88 311.42 930.86 ;
     RECT  311.14 1425.84 312.1 1430.66 ;
     RECT  311.42 923.1 312.38 930.86 ;
     RECT  312.1 1425.84 313.54 1426.04 ;
     RECT  306.82 1368.285 313.955 1369.76 ;
     RECT  310.18 1440.12 314.02 1479.76 ;
     RECT  310.46 941.58 314.3 1350.875 ;
     RECT  312.38 921.84 314.78 930.86 ;
     RECT  314.3 940.74 314.78 1350.875 ;
     RECT  313.955 1368.3 314.98 1369.76 ;
     RECT  314.78 921.84 315.26 1350.875 ;
     RECT  311.19 215.36 316.81 878.32 ;
     RECT  311.19 1577 316.81 1583.92 ;
     RECT  315.26 921.84 319.1 1355.06 ;
     RECT  319.1 918.9 322.46 1355.06 ;
     RECT  322.46 918.9 322.94 1356.74 ;
     RECT  314.02 1440.12 323.42 1470.98 ;
     RECT  314.02 1479.56 323.42 1479.76 ;
     RECT  323.42 1439.7 323.62 1479.76 ;
     RECT  322.94 918.9 323.9 1357.58 ;
     RECT  314.98 1368.3 323.9 1368.5 ;
     RECT  316.81 1577 327.74 1578.04 ;
     RECT  323.9 918.9 332.455 1368.5 ;
     RECT  323.62 1447.26 333.02 1479.76 ;
     RECT  332.455 915.96 333.235 1368.5 ;
     RECT  333.235 915.12 336.745 1368.5 ;
     RECT  336.745 915.12 337.24 1376.075 ;
     RECT  337.24 915.12 337.34 1376.91 ;
     RECT  337.34 915.12 338.24 1379.84 ;
     RECT  316.81 615.62 338.78 616.66 ;
     RECT  338.78 1430.04 339.26 1434.02 ;
     RECT  338.78 1392.24 339.68 1392.44 ;
     RECT  339.26 1430.04 339.68 1436.96 ;
     RECT  338.24 915.12 339.74 1380.85 ;
     RECT  339.68 1391.23 339.74 1392.44 ;
     RECT  339.68 1429.03 340.16 1436.96 ;
     RECT  340.16 1429.03 341.6 1436.995 ;
     RECT  333.02 1445.58 341.6 1479.76 ;
     RECT  339.74 915.12 343.58 1392.44 ;
     RECT  341.6 1429.03 344.06 1479.76 ;
     RECT  343.58 915.12 345.5 1394.54 ;
     RECT  345.5 915.12 346.94 1399.16 ;
     RECT  338.78 615.62 347.42 619.6 ;
     RECT  346.94 915.12 347.42 1400.84 ;
     RECT  347.42 914.28 347.9 1400.84 ;
     RECT  344.06 1425.84 348.86 1479.76 ;
     RECT  348.86 1417.86 353.66 1479.76 ;
     RECT  347.9 906.72 354.985 1400.84 ;
     RECT  353.66 1409.88 354.985 1479.76 ;
     RECT  293 -70 363 180 ;
     RECT  293 1620 363 1870 ;
     RECT  354.985 906.72 364.42 1479.76 ;
     RECT  316.81 388.4 379.19 563.74 ;
     RECT  316.81 588.74 379.19 588.94 ;
     RECT  347.42 614.78 379.19 619.6 ;
     RECT  316.81 629.9 379.19 630.1 ;
     RECT  316.81 651.32 379.19 651.52 ;
     RECT  316.81 673.16 379.19 673.36 ;
     RECT  316.81 684.5 379.19 837.58 ;
     RECT  316.81 857.54 379.19 878.32 ;
     RECT  327.74 1577 379.19 1578.46 ;
     RECT  364.42 907.14 380.26 1479.76 ;
     RECT  363 0 381 180 ;
     RECT  363 1620 381 1800 ;
     RECT  379.19 219.14 384.81 878.32 ;
     RECT  379.19 1577 384.81 1580.14 ;
     RECT  380.26 907.56 395.84 1479.76 ;
     RECT  397.82 219.98 402.14 221.44 ;
     RECT  395.84 907.39 403.285 1479.76 ;
     RECT  402.14 217.46 403.58 221.44 ;
     RECT  403.58 217.46 405.22 225.22 ;
     RECT  405.22 217.46 407.14 222.28 ;
     RECT  384.81 388.4 407.9 563.74 ;
     RECT  407.14 217.46 408.1 217.66 ;
     RECT  384.81 629.9 409.34 630.1 ;
     RECT  405.5 639.14 409.34 639.34 ;
     RECT  403.285 908.4 412.435 1479.76 ;
     RECT  412.435 907.56 414.34 1479.76 ;
     RECT  381 1620 417.5 1870 ;
     RECT  417.5 1619.42 417.7 1870 ;
     RECT  414.34 907.56 421.29 1478.96 ;
     RECT  407.9 388.4 426.14 565.84 ;
     RECT  421.29 907.98 430.46 1478.96 ;
     RECT  430.46 906.3 433.82 1478.96 ;
     RECT  384.81 673.16 437.18 673.36 ;
     RECT  384.81 1577 439.1 1578.46 ;
     RECT  433.82 906.3 440.74 1479.38 ;
     RECT  384.81 857.54 441.02 878.32 ;
     RECT  440.74 906.3 442.18 1478.96 ;
     RECT  442.18 906.3 443.14 1478.12 ;
     RECT  441.02 857.54 443.42 881.3 ;
     RECT  443.14 906.3 445.82 1448.3 ;
     RECT  443.14 1459.27 448.405 1478.12 ;
     RECT  448.405 1460.7 449.86 1478.12 ;
     RECT  381 -70 451 180 ;
     RECT  417.7 1620 451 1870 ;
     RECT  449.86 1460.7 451.78 1471.4 ;
     RECT  409.34 629.9 454.94 639.34 ;
     RECT  445.82 898.32 455.9 1448.3 ;
     RECT  454.94 629.9 460.22 642.7 ;
     RECT  384.81 651.32 460.22 651.52 ;
     RECT  455.9 898.32 460.42 1452.08 ;
     RECT  460.42 898.32 460.9 1447.88 ;
     RECT  460.22 629.9 463.58 651.52 ;
     RECT  460.9 898.32 467.14 1447.46 ;
     RECT  451 0 469 180 ;
     RECT  451 1620 469 1800 ;
     RECT  443.42 857.54 470.3 882.14 ;
     RECT  467.14 1435.92 470.98 1447.46 ;
     RECT  384.81 614.78 473.18 619.6 ;
     RECT  467.14 898.32 473.86 1426.21 ;
     RECT  473.86 1364.1 474.325 1426.21 ;
     RECT  474.325 1364.1 474.82 1425.62 ;
     RECT  470.98 1435.92 475.715 1441.595 ;
     RECT  475.715 1435.92 476.165 1440.76 ;
     RECT  474.82 1364.1 476.26 1425.2 ;
     RECT  476.165 1435.92 476.74 1440.74 ;
     RECT  451.78 1471.2 476.74 1471.4 ;
     RECT  476.74 1435.92 477.22 1436.12 ;
     RECT  473.86 898.32 477.685 1353.8 ;
     RECT  476.26 1424.58 477.7 1425.2 ;
     RECT  439.1 1577 478.46 1582.24 ;
     RECT  477.685 898.32 481.06 1350.44 ;
     RECT  473.18 608.9 481.34 619.6 ;
     RECT  463.58 629.9 481.34 654.46 ;
     RECT  437.18 673.16 481.34 674.2 ;
     RECT  384.81 682.82 481.34 837.58 ;
     RECT  469 -70 485.42 180 ;
     RECT  485.42 -70 485.86 180.7 ;
     RECT  481.06 1250.7 486.14 1350.44 ;
     RECT  476.26 1364.1 486.14 1411.09 ;
     RECT  486.14 1250.7 488.54 1419.78 ;
     RECT  486.14 1429.24 488.54 1431.12 ;
     RECT  486.14 1442.26 488.54 1442.46 ;
     RECT  481.06 898.32 489.515 1242.12 ;
     RECT  488.54 1250.7 489.515 1431.12 ;
     RECT  488.54 1440.16 489.515 1447.5 ;
     RECT  478.46 1577 489.7 1582.66 ;
     RECT  481.34 608.9 489.98 654.46 ;
     RECT  489.515 898.32 491.515 1447.5 ;
     RECT  491.515 898.32 493.82 1447.51 ;
     RECT  490.94 1464.94 495.74 1465.14 ;
     RECT  470.3 857.54 496.42 884.66 ;
     RECT  493.82 898.32 497.18 1455.9 ;
     RECT  495.74 1464.94 497.18 1468.92 ;
     RECT  497.18 898.32 499.115 1468.92 ;
     RECT  499.115 898.32 502.18 1469.76 ;
     RECT  502.18 1169.26 502.335 1469.76 ;
     RECT  502.335 1169.26 502.94 1473.54 ;
     RECT  489.98 608.9 504.38 662.02 ;
     RECT  481.34 673.16 504.38 837.58 ;
     RECT  469 1620 505.34 1870 ;
     RECT  505.34 1619.42 506.5 1870 ;
     RECT  502.18 898.32 513.02 1157.24 ;
     RECT  485.66 223.34 515.19 223.54 ;
     RECT  426.14 388.4 515.19 567.52 ;
     RECT  384.81 588.74 515.19 588.94 ;
     RECT  426.62 600.08 515.19 600.28 ;
     RECT  504.38 608.9 515.19 837.58 ;
     RECT  496.42 857.54 515.19 882.14 ;
     RECT  489.7 1577 515.19 1582.24 ;
     RECT  502.94 1169.26 518.3 1478.16 ;
     RECT  515.19 215.36 520.81 882.14 ;
     RECT  515.19 1577 520.81 1583.92 ;
     RECT  513.02 891.18 521.66 1157.24 ;
     RECT  518.3 1169.26 521.66 1481.1 ;
     RECT  521.66 891.18 525.98 1481.1 ;
     RECT  525.98 891.18 527.62 1482.36 ;
     RECT  527.62 1152.46 530.02 1482.36 ;
     RECT  530.02 1152.46 537.22 1481.94 ;
     RECT  527.62 891.18 537.7 1143.38 ;
     RECT  537.22 1152.46 538.29 1481.1 ;
     RECT  485.86 -70 539 180 ;
     RECT  506.5 1620 539 1870 ;
     RECT  538.29 1152.46 545.86 1480.26 ;
     RECT  545.86 1152.46 550.66 1478.58 ;
     RECT  550.66 1152.46 551.2 1477.355 ;
     RECT  539 0 557 180 ;
     RECT  539 1620 557 1800 ;
     RECT  551.2 1152.46 561.02 1477.32 ;
     RECT  561.02 1152.04 561.5 1477.32 ;
     RECT  561.5 1152.04 567.26 1477.74 ;
     RECT  557 -70 570.38 180 ;
     RECT  567.26 1152.04 570.635 1480.26 ;
     RECT  570.38 -70 570.82 180.7 ;
     RECT  520.81 223.34 573.5 223.54 ;
     RECT  570.635 1152.04 580.7 1481.69 ;
     RECT  580.7 1152.04 581.66 1484.88 ;
     RECT  573.5 223.34 583.19 224.38 ;
     RECT  520.81 388.4 583.19 567.52 ;
     RECT  520.81 588.74 583.19 588.94 ;
     RECT  520.81 600.08 583.19 600.28 ;
     RECT  520.81 608.9 583.19 837.58 ;
     RECT  520.81 857.54 583.19 882.14 ;
     RECT  581.66 1152.04 583.58 1485.3 ;
     RECT  232.22 1493.84 583.58 1494.04 ;
     RECT  583.58 1152.04 586.46 1494.04 ;
     RECT  583.19 219.14 588.81 882.14 ;
     RECT  557 1620 593.18 1870 ;
     RECT  586.46 1151.62 593.38 1494.04 ;
     RECT  593.18 1619.42 593.38 1870 ;
     RECT  593.38 1151.62 595.3 1485.3 ;
     RECT  588.81 600.08 597.7 842.2 ;
     RECT  588.81 388.4 605.66 567.52 ;
     RECT  605.66 388.4 606.14 569.62 ;
     RECT  606.14 388.4 606.62 570.04 ;
     RECT  606.62 388.4 608.06 570.88 ;
     RECT  595.3 1151.62 609.5 1482.36 ;
     RECT  608.06 388.4 610.46 577.18 ;
     RECT  610.46 388.4 611.36 579.7 ;
     RECT  588.81 588.74 611.36 588.94 ;
     RECT  570.82 -70 611.9 180 ;
     RECT  611.9 -70 612.1 180.7 ;
     RECT  597.7 608.06 612.295 842.2 ;
     RECT  612.295 606.8 612.38 842.2 ;
     RECT  612.38 603.86 613.34 842.2 ;
     RECT  537.7 891.18 614.02 1138.76 ;
     RECT  611.36 388.4 614.3 588.94 ;
     RECT  613.34 602.6 614.3 842.2 ;
     RECT  609.5 1149.52 614.98 1482.36 ;
     RECT  614.3 388.4 619.3 842.2 ;
     RECT  588.81 857.54 619.3 882.14 ;
     RECT  619.3 857.96 623.42 882.14 ;
     RECT  614.98 1149.52 623.9 1481.1 ;
     RECT  623.9 1149.52 625.34 1481.52 ;
     RECT  612.1 -70 627 180 ;
     RECT  593.38 1620 627 1870 ;
     RECT  625.34 1148.26 636.86 1481.52 ;
     RECT  614.02 898.32 639.26 1138.76 ;
     RECT  636.86 1148.26 639.26 1481.94 ;
     RECT  520.81 1577 640.9 1582.24 ;
     RECT  639.26 898.32 641.38 1481.94 ;
     RECT  641.38 898.32 643.3 1481.1 ;
     RECT  627 0 645 180 ;
     RECT  627 1620 645 1800 ;
     RECT  619.3 388.4 647.42 839.68 ;
     RECT  623.42 857.96 652.615 887.6 ;
     RECT  647.42 388.4 652.7 842.2 ;
     RECT  652.615 851.66 652.7 887.6 ;
     RECT  652.7 388.4 653.86 887.6 ;
     RECT  643.3 898.32 666.14 1478.16 ;
     RECT  588.81 223.34 666.62 224.38 ;
     RECT  233.66 1558.52 666.82 1565.86 ;
     RECT  653.86 887.4 668.74 887.6 ;
     RECT  666.62 220.82 672.58 224.38 ;
     RECT  666.14 898.32 673.06 1481.52 ;
     RECT  673.06 898.32 674.98 1480.68 ;
     RECT  653.86 388.4 676.22 878.32 ;
     RECT  645 1620 677.66 1870 ;
     RECT  677.66 1619.42 678.82 1870 ;
     RECT  674.98 898.32 681.7 1478.16 ;
     RECT  676.22 388.4 685.82 886.76 ;
     RECT  681.7 898.32 685.82 1475.22 ;
     RECT  640.9 1577 691.3 1581.82 ;
     RECT  685.82 388.4 692.26 1475.22 ;
     RECT  692.26 903.36 693.7 1473.54 ;
     RECT  693.7 903.36 701.38 1472.28 ;
     RECT  692.26 388.4 702.34 894.74 ;
     RECT  702.34 388.4 706.66 886.76 ;
     RECT  701.38 1152.46 708.58 1472.28 ;
     RECT  701.38 903.36 714.34 1139.22 ;
     RECT  645 -70 715 180 ;
     RECT  678.82 1620 715 1870 ;
     RECT  672.58 223.34 719.19 224.38 ;
     RECT  706.66 388.4 719.19 879.16 ;
     RECT  691.3 1577 719.19 1580.98 ;
     RECT  708.58 1152.46 721.82 1471.02 ;
     RECT  714.34 903.36 724.22 1138.8 ;
     RECT  719.19 215.36 724.81 879.16 ;
     RECT  719.19 1577 724.81 1583.92 ;
     RECT  721.82 1152.46 726.635 1473.96 ;
     RECT  724.81 388.4 729.7 879.16 ;
     RECT  715 0 733 180 ;
     RECT  715 1620 733 1800 ;
     RECT  726.635 1152.46 734.08 1474.13 ;
     RECT  734.08 1152.46 734.3 1473.12 ;
     RECT  729.7 388.4 734.5 878.32 ;
     RECT  734.3 1152.04 735.46 1473.12 ;
     RECT  724.22 903.36 738.82 1143 ;
     RECT  734.5 605.96 741.5 878.32 ;
     RECT  724.81 1577 741.5 1580.98 ;
     RECT  741.5 605.96 743.42 878.74 ;
     RECT  738.82 904.62 745.34 1143 ;
     RECT  735.46 1152.04 745.82 1471.44 ;
     RECT  734.5 388.4 748.7 597.34 ;
     RECT  743.42 605.96 748.7 879.16 ;
     RECT  733 -70 749.42 180 ;
     RECT  724.81 223.34 749.66 224.38 ;
     RECT  745.82 1152.04 749.66 1473.96 ;
     RECT  749.42 -70 749.86 180.7 ;
     RECT  745.34 904.62 753.22 1143.42 ;
     RECT  749.66 219.98 755.62 224.38 ;
     RECT  753.22 904.62 765.5 1138.8 ;
     RECT  748.7 388.4 767.9 879.16 ;
     RECT  749.66 1152.04 775.3 1479.76 ;
     RECT  775.3 1153.3 776.26 1479.76 ;
     RECT  776.26 1153.72 780.1 1479.76 ;
     RECT  780.1 1154.14 786.62 1479.76 ;
     RECT  765.5 903.78 786.82 1138.8 ;
     RECT  755.62 223.34 787.19 224.38 ;
     RECT  767.9 388.4 787.19 880.42 ;
     RECT  786.82 904.2 792.1 1138.8 ;
     RECT  792.1 904.62 792.58 1138.8 ;
     RECT  787.19 219.14 792.81 880.42 ;
     RECT  786.62 1154.14 794.08 1480.18 ;
     RECT  749.86 -70 803 180 ;
     RECT  733 1620 803 1870 ;
     RECT  794.08 1154.14 805.06 1470.6 ;
     RECT  805.06 1154.56 805.54 1470.6 ;
     RECT  792.81 388.4 805.82 880.42 ;
     RECT  792.58 906.3 806.5 1138.8 ;
     RECT  805.54 1154.56 806.98 1470.18 ;
     RECT  806.98 1154.56 808.9 1469.34 ;
     RECT  806.5 906.3 817.78 1137.96 ;
     RECT  817.78 906.3 820.42 1064 ;
     RECT  808.9 1154.56 820.48 1466.57 ;
     RECT  803 0 821 180 ;
     RECT  803 1620 821 1800 ;
     RECT  820.48 1154.56 821.38 1465.56 ;
     RECT  805.82 388.4 822.82 887.6 ;
     RECT  821.38 1154.56 822.82 1463.88 ;
     RECT  820.42 907.98 824.74 1064 ;
     RECT  817.78 1074.3 824.74 1137.96 ;
     RECT  822.82 1157.08 826.18 1463.88 ;
     RECT  824.74 1082.28 826.66 1127 ;
     RECT  826.66 1082.7 827.14 1127 ;
     RECT  827.14 1082.7 827.62 1123.22 ;
     RECT  827.62 1082.7 828.1 1122.38 ;
     RECT  822.82 388.4 829.06 885.5 ;
     RECT  828.1 1083.12 829.54 1122.38 ;
     RECT  826.18 1160.86 830.02 1463.88 ;
     RECT  829.06 614.78 831.26 885.5 ;
     RECT  829.54 1083.12 831.46 1121.54 ;
     RECT  831.46 1084.38 831.94 1121.54 ;
     RECT  831.94 1084.38 832.18 1116.92 ;
     RECT  832.18 1084.38 832.66 1116.08 ;
     RECT  832.66 1089.42 832.9 1116.08 ;
     RECT  832.9 1089.42 833.38 1114.82 ;
     RECT  833.38 1090.26 833.62 1114.82 ;
     RECT  824.74 1137.76 833.86 1137.96 ;
     RECT  833.62 1090.26 834.34 1107.68 ;
     RECT  821 -70 834.38 180 ;
     RECT  831.26 614.78 834.62 885.92 ;
     RECT  794.08 1479.56 834.62 1480.18 ;
     RECT  834.38 -70 834.82 180.7 ;
     RECT  834.34 1092.78 834.82 1107.68 ;
     RECT  824.74 907.98 836.245 1063.33 ;
     RECT  834.82 1092.78 836.26 1107.26 ;
     RECT  836.26 1092.78 837.22 1105.16 ;
     RECT  792.81 223.34 837.5 224.38 ;
     RECT  837.22 1093.62 837.7 1105.16 ;
     RECT  837.7 1093.62 838.66 1096.76 ;
     RECT  838.66 1093.62 839.14 1095.08 ;
     RECT  839.14 1093.62 839.38 1093.82 ;
     RECT  836.245 907.98 839.62 1061.9 ;
     RECT  834.62 614.78 840.1 886.34 ;
     RECT  830.02 1161.7 841.06 1463.88 ;
     RECT  841.06 1161.7 841.54 1161.9 ;
     RECT  837.5 219.98 843.94 224.38 ;
     RECT  841.06 1175.14 844.7 1463.88 ;
     RECT  834.62 1472.42 844.7 1480.18 ;
     RECT  839.62 907.98 844.9 1060.22 ;
     RECT  840.1 614.78 846.82 885.92 ;
     RECT  844.9 907.98 847.78 1058.96 ;
     RECT  829.06 388.4 849.34 604.48 ;
     RECT  849.34 388.4 849.5 606.16 ;
     RECT  846.82 614.78 849.5 880.42 ;
     RECT  847.78 915.12 851.125 1058.96 ;
     RECT  851.125 915.12 854.5 1058.12 ;
     RECT  741.5 1577 855.94 1582.24 ;
     RECT  844.7 1175.14 856.9 1480.18 ;
     RECT  854.5 915.12 857.86 1057.7 ;
     RECT  857.86 915.12 858.34 1054.34 ;
     RECT  858.34 915.12 858.82 1048.21 ;
     RECT  858.82 915.96 862.645 1048.21 ;
     RECT  856.9 1175.14 862.66 1462.62 ;
     RECT  862.645 915.96 865.06 1047.2 ;
     RECT  862.66 1175.14 867.46 1458.42 ;
     RECT  867.46 1175.14 868.9 1451.45 ;
     RECT  868.9 1189.84 869.38 1451.45 ;
     RECT  869.38 1192.78 869.86 1451.45 ;
     RECT  869.86 1192.78 870.82 1440.36 ;
     RECT  869.86 1450.24 870.88 1451.45 ;
     RECT  870.88 1450.24 871.78 1450.44 ;
     RECT  865.06 918.9 871.945 1047.2 ;
     RECT  870.82 1193.62 872.74 1440.36 ;
     RECT  872.74 1197.82 873.22 1440.36 ;
     RECT  834.82 -70 875.9 180 ;
     RECT  821 1620 875.9 1870 ;
     RECT  875.9 -70 876.1 180.7 ;
     RECT  871.945 918.9 876.1 1048.475 ;
     RECT  875.9 1619.42 876.1 1870 ;
     RECT  876.1 918.9 876.58 1036.7 ;
     RECT  876.58 918.9 878.5 919.1 ;
     RECT  873.22 1197.82 878.98 1432.72 ;
     RECT  876.1 1047 879.395 1048.475 ;
     RECT  878.98 1424.62 879.46 1432.72 ;
     RECT  879.395 1047 879.845 1047.64 ;
     RECT  876.58 931.92 880.42 1036.7 ;
     RECT  879.845 1047 880.42 1047.62 ;
     RECT  878.98 1197.82 880.42 1416 ;
     RECT  849.5 388.4 880.7 880.42 ;
     RECT  880.42 1348.43 880.9 1416 ;
     RECT  880.7 388.4 881.18 885.46 ;
     RECT  880.42 935.28 881.38 1036.7 ;
     RECT  880.9 1406.56 881.38 1416 ;
     RECT  880.42 1197.82 881.86 1338.05 ;
     RECT  880.9 1348.43 881.86 1397.52 ;
     RECT  881.38 1406.56 881.86 1412.22 ;
     RECT  881.38 942.84 882.34 1036.7 ;
     RECT  881.86 1197.82 882.34 1219.86 ;
     RECT  881.86 1242.34 882.34 1338.05 ;
     RECT  881.86 1372.12 882.34 1387.44 ;
     RECT  881.86 1348.43 882.4 1360.73 ;
     RECT  882.34 1197.82 882.62 1217.09 ;
     RECT  882.34 959.64 882.82 1036.7 ;
     RECT  882.34 1242.34 882.82 1326.155 ;
     RECT  881.86 1406.56 882.88 1409.315 ;
     RECT  881.18 388.4 883.1 885.88 ;
     RECT  882.82 1242.34 883.3 1269.42 ;
     RECT  882.34 1378 883.3 1387.44 ;
     RECT  882.82 1288.12 883.36 1326.155 ;
     RECT  882.34 1336.84 883.36 1338.05 ;
     RECT  882.4 1348.43 883.36 1356.78 ;
     RECT  882.62 1142.72 883.58 1142.92 ;
     RECT  882.34 942.84 883.78 948.5 ;
     RECT  882.88 1406.56 883.78 1409.28 ;
     RECT  883.3 1242.34 883.84 1254.72 ;
     RECT  883.36 1288.12 883.84 1323.6 ;
     RECT  883.3 1386.23 883.84 1387.44 ;
     RECT  882.62 1194.38 884.06 1217.09 ;
     RECT  883.78 948.3 884.26 948.5 ;
     RECT  884.06 1190.6 884.26 1217.09 ;
     RECT  883.84 1254.1 884.26 1254.72 ;
     RECT  883.84 1288.12 884.26 1291.68 ;
     RECT  883.84 1315.84 884.26 1323.6 ;
     RECT  883.36 1336.84 884.26 1337.04 ;
     RECT  883.36 1349.44 884.26 1356.78 ;
     RECT  883.84 1242.34 884.74 1244.14 ;
     RECT  884.26 1288.12 884.74 1288.32 ;
     RECT  883.84 1300.72 884.74 1300.92 ;
     RECT  884.26 1315.84 884.74 1323.52 ;
     RECT  883.84 1387.24 884.74 1387.44 ;
     RECT  883.1 1156.16 885.5 1156.36 ;
     RECT  882.82 959.64 886.18 1035.44 ;
     RECT  855.94 1577 889.06 1578.04 ;
     RECT  886.18 959.64 890.02 1033.76 ;
     RECT  889.06 1577.42 890.02 1578.04 ;
     RECT  876.1 -70 891 180 ;
     RECT  876.1 1620 891 1870 ;
     RECT  884.26 1214.12 891.26 1217.09 ;
     RECT  884.26 1190.6 892.22 1196.68 ;
     RECT  883.1 388.4 892.7 887.98 ;
     RECT  892.7 388.4 892.9 891.34 ;
     RECT  883.58 1136.42 894.14 1142.92 ;
     RECT  885.5 1156.16 894.62 1164.76 ;
     RECT  892.22 1182.62 894.62 1196.68 ;
     RECT  891.26 1214.12 895.58 1218.1 ;
     RECT  893.18 904.58 896.54 904.78 ;
     RECT  894.62 1156.16 896.54 1166.86 ;
     RECT  894.62 1182.2 896.54 1196.68 ;
     RECT  884.26 1352.3 896.54 1352.5 ;
     RECT  896.54 1344.32 897.02 1352.5 ;
     RECT  890.02 1577.84 897.035 1578.04 ;
     RECT  892.9 648.38 897.5 891.34 ;
     RECT  896.54 904.58 897.5 905.2 ;
     RECT  895.58 923.9 897.5 924.1 ;
     RECT  896.06 932.72 897.5 932.92 ;
     RECT  890.02 959.64 897.5 1029.98 ;
     RECT  894.14 1136.42 897.5 1144.6 ;
     RECT  897.035 1577.84 897.865 1580.14 ;
     RECT  897.5 648.38 897.98 905.2 ;
     RECT  891.74 914.24 897.98 914.44 ;
     RECT  897.5 923.9 897.98 934.6 ;
     RECT  897.5 952.88 897.98 1029.98 ;
     RECT  897.5 1129.28 897.98 1144.6 ;
     RECT  896.54 1156.16 897.98 1196.68 ;
     RECT  895.58 1209.92 897.98 1218.1 ;
     RECT  897.865 1577.84 898.36 1581.415 ;
     RECT  897.02 1260.74 900.38 1260.94 ;
     RECT  897.98 648.38 900.775 1029.98 ;
     RECT  879.46 1432.52 901.035 1432.72 ;
     RECT  856.9 1472.42 901.035 1480.18 ;
     RECT  593.38 1493.84 901.035 1494.04 ;
     RECT  222.62 1544.24 901.035 1544.44 ;
     RECT  666.82 1565.66 901.035 1565.86 ;
     RECT  898.36 1577.84 901.035 1582.25 ;
     RECT  900.775 648.38 902.3 1030.78 ;
     RECT  902.3 648.38 902.78 1034.14 ;
     RECT  884.74 1243.94 902.78 1244.14 ;
     RECT  901.035 1372.04 902.965 1583.92 ;
     RECT  902.3 1081.4 903.26 1083.7 ;
     RECT  902.78 1093.16 903.26 1094.2 ;
     RECT  900.38 1260.74 903.26 1262.62 ;
     RECT  902.965 1565.66 903.46 1565.86 ;
     RECT  902.78 1239.32 903.74 1244.14 ;
     RECT  902.965 1577.84 903.94 1582.25 ;
     RECT  899.9 1227.56 904.22 1227.76 ;
     RECT  903.74 1237.22 904.22 1244.14 ;
     RECT  902.965 1408.16 904.42 1544.44 ;
     RECT  903.26 1260.74 904.7 1263.88 ;
     RECT  903.74 1274.18 904.7 1274.38 ;
     RECT  904.22 1045.28 905.18 1048 ;
     RECT  903.26 1056.62 905.18 1056.82 ;
     RECT  896.06 1307.78 905.18 1307.98 ;
     RECT  884.74 1323.32 905.18 1323.52 ;
     RECT  897.02 1336.76 905.18 1352.5 ;
     RECT  903.94 1581.185 905.315 1582.25 ;
     RECT  903.26 1081.4 905.66 1094.2 ;
     RECT  902.3 1112.9 905.66 1113.1 ;
     RECT  897.98 1129.28 905.66 1218.1 ;
     RECT  902.965 1372.04 905.66 1378.12 ;
     RECT  905.315 1581.2 905.765 1582.25 ;
     RECT  905.095 1070.9 905.875 1071.1 ;
     RECT  905.18 1044.86 906.62 1056.82 ;
     RECT  905.66 1112.9 906.62 1218.1 ;
     RECT  904.22 1227.56 906.62 1251.7 ;
     RECT  905.765 1581.2 906.82 1581.4 ;
     RECT  906.62 1044.86 906.94 1060.6 ;
     RECT  905.875 1070.9 906.94 1071.94 ;
     RECT  902.78 648.38 906.975 1035.4 ;
     RECT  906.94 1044.86 906.975 1071.94 ;
     RECT  905.66 1080.98 907.04 1094.2 ;
     RECT  892.9 388.4 907.1 638.5 ;
     RECT  906.975 648.38 907.1 1071.94 ;
     RECT  895.1 1293.08 907.1 1293.28 ;
     RECT  905.18 1307.78 907.1 1309.66 ;
     RECT  905.66 1371.2 907.1 1378.12 ;
     RECT  907.04 1080.98 907.58 1098.015 ;
     RECT  906.62 1112.9 907.58 1251.7 ;
     RECT  904.7 1260.74 907.58 1274.38 ;
     RECT  907.1 388.4 908 1071.94 ;
     RECT  907.58 1080.56 908 1098.015 ;
     RECT  908 388.4 908.06 1098.015 ;
     RECT  907.58 1112.9 908.06 1274.38 ;
     RECT  907.1 1283.42 908.06 1283.62 ;
     RECT  907.1 1293.08 908.06 1309.66 ;
     RECT  905.18 1323.32 908.06 1352.5 ;
     RECT  907.1 1363.64 908.06 1378.12 ;
     RECT  891 0 909 180 ;
     RECT  891 1620 909 1800 ;
     RECT  908.06 1283 909.5 1283.62 ;
     RECT  908.06 1293.08 909.5 1378.12 ;
     RECT  908.06 1108.7 910.7 1274.38 ;
     RECT  909.5 1283 910.7 1378.12 ;
     RECT  910.7 1108.7 914.3 1378.12 ;
     RECT  904.42 1408.16 914.78 1543.18 ;
     RECT  911.9 1554.32 914.78 1554.52 ;
     RECT  908.06 388.4 915.26 1098.4 ;
     RECT  914.3 1107.02 915.26 1378.12 ;
     RECT  914.78 1407.74 915.99 1557.04 ;
     RECT  915.99 1399.075 918.155 1557.04 ;
     RECT  918.155 1399.075 918.62 1558.47 ;
     RECT  918.62 1399.075 918.8 1561.66 ;
     RECT  918.8 1398.58 919.1 1561.66 ;
     RECT  915.26 388.4 919.58 1378.12 ;
     RECT  912.38 1386.74 919.58 1386.94 ;
     RECT  919.58 388.4 921.02 1386.94 ;
     RECT  919.1 1396.4 921.02 1561.66 ;
     RECT  843.94 223.34 923.19 224.38 ;
     RECT  921.02 388.4 923.19 1561.66 ;
     RECT  923.19 215.36 924.38 1561.66 ;
     RECT  924.38 215.36 927.26 1562.08 ;
     RECT  927.26 215.36 928.81 1569.64 ;
     RECT  923.19 1583.72 928.81 1583.92 ;
     RECT  928.81 388.4 935.14 1569.64 ;
     RECT  935.14 408.98 938.5 1569.64 ;
     RECT  938.5 409.4 939.94 1569.64 ;
     RECT  939.94 409.4 942.82 1568.38 ;
     RECT  935.14 388.4 950.02 395.74 ;
     RECT  942.82 409.82 953.86 1562.5 ;
     RECT  953.86 409.82 956.26 1559.14 ;
     RECT  956.26 658.46 956.74 1559.14 ;
     RECT  956.26 409.82 957.7 649 ;
     RECT  956.54 1568.85 959.915 1572.16 ;
     RECT  957.7 409.82 960.58 648.58 ;
     RECT  960.58 410.24 964.42 648.58 ;
     RECT  964.42 416.12 966.62 648.58 ;
     RECT  956.74 660.98 966.62 1559.14 ;
     RECT  966.62 416.12 968.06 1559.14 ;
     RECT  959.915 1568.85 968.06 1573.59 ;
     RECT  968.06 416.12 969.02 1573.59 ;
     RECT  969.02 416.12 969.7 1577.62 ;
     RECT  969.7 416.96 971.42 1577.62 ;
     RECT  909 -70 979 180 ;
     RECT  909 1620 979 1870 ;
     RECT  971.42 416.96 982.66 1578.04 ;
     RECT  928.81 223.34 991.19 224.38 ;
     RECT  950.02 388.4 991.19 392.8 ;
     RECT  982.66 416.96 991.19 1577.62 ;
     RECT  991.19 219.14 996.81 1580.14 ;
     RECT  979 0 997 180 ;
     RECT  979 1620 997 1800 ;
     RECT  996.81 423.68 998.02 1577.62 ;
     RECT  998.02 666.86 1002.82 1577.62 ;
     RECT  996.81 388.4 1005.22 392.8 ;
     RECT  1002.82 669.8 1005.5 1577.62 ;
     RECT  998.02 423.68 1007.42 656.98 ;
     RECT  1007.42 423.68 1009.555 659.5 ;
     RECT  1009.555 423.26 1011.485 659.5 ;
     RECT  1011.485 423.68 1012.42 423.88 ;
     RECT  1011.485 519.44 1012.42 659.5 ;
     RECT  1005.5 669.8 1012.7 1581.82 ;
     RECT  1012.42 519.86 1013.18 659.5 ;
     RECT  1012.7 669.8 1013.18 1583.08 ;
     RECT  997 -70 1013.42 180 ;
     RECT  996.81 223.34 1013.66 224.38 ;
     RECT  1013.42 -70 1013.86 180.7 ;
     RECT  1005.22 392.6 1013.86 392.8 ;
     RECT  1013.18 519.86 1015.765 1583.08 ;
     RECT  1015.765 520.7 1019.14 1583.08 ;
     RECT  1013.66 219.98 1020.58 224.38 ;
     RECT  1019.14 524.48 1021.54 1583.08 ;
     RECT  1021.54 527.42 1026.805 1583.08 ;
     RECT  1026.805 530.61 1030.165 1583.08 ;
     RECT  1030.165 532.04 1031.125 1583.08 ;
     RECT  1031.125 532.04 1033.54 533.92 ;
     RECT  1033.54 533.72 1034.5 533.92 ;
     RECT  1031.125 543.38 1034.5 1583.08 ;
     RECT  1034.5 545.9 1043.9 1583.08 ;
     RECT  1020.58 223.34 1044.1 224.38 ;
     RECT  1043.9 545.9 1049.86 1583.5 ;
     RECT  1049.86 545.9 1052.74 1583.08 ;
     RECT  1044.1 223.76 1053.22 224.38 ;
     RECT  1052.74 545.9 1053.22 1050.1 ;
     RECT  1052.74 1060.4 1055.62 1583.08 ;
     RECT  1053.22 546.32 1056.1 1050.1 ;
     RECT  1056.1 547.16 1060.9 1050.1 ;
     RECT  1060.9 655.52 1063.58 1050.1 ;
     RECT  1055.62 1060.4 1063.58 1582.66 ;
     RECT  1063.58 655.52 1065.22 1582.66 ;
     RECT  1060.9 547.16 1066.22 646.9 ;
     RECT  1013.86 -70 1067 180 ;
     RECT  997 1620 1067 1870 ;
     RECT  1066.22 546.32 1067.305 646.9 ;
     RECT  1067.305 545.465 1069.82 646.9 ;
     RECT  1065.22 655.52 1069.82 1582.24 ;
     RECT  1069.82 545.465 1073.62 1582.24 ;
     RECT  1073.62 545.465 1074.755 1056.4 ;
     RECT  1074.755 546.3 1075.205 1056.4 ;
     RECT  1053.22 223.76 1078.66 223.96 ;
     RECT  1075.205 546.32 1080.58 1056.4 ;
     RECT  1080.58 659.13 1082.005 1056.4 ;
     RECT  1073.62 1066.28 1082.5 1582.24 ;
     RECT  1082.005 660.14 1082.78 1056.4 ;
     RECT  1082.5 1066.28 1082.78 1566.03 ;
     RECT  1082.78 660.14 1084.42 1566.03 ;
     RECT  1084.42 660.56 1084.9 1566.03 ;
     RECT  1067 0 1085 180 ;
     RECT  1067 1620 1085 1800 ;
     RECT  1084.9 660.56 1085.38 1549.48 ;
     RECT  1080.58 546.32 1085.42 648.58 ;
     RECT  1085.38 662.24 1085.94 1549.48 ;
     RECT  1085.94 662.24 1086.42 1527.22 ;
     RECT  1084.9 1564.82 1086.88 1566.03 ;
     RECT  1086.42 662.24 1087.75 1524.62 ;
     RECT  1086.88 1564.82 1087.78 1565.02 ;
     RECT  1085.42 545.9 1090.94 648.58 ;
     RECT  1085.94 1539.2 1091.14 1549.48 ;
     RECT  1090.94 542.12 1092.38 648.58 ;
     RECT  1091.14 1539.2 1093.06 1549.06 ;
     RECT  1092.38 540.44 1093.28 651.94 ;
     RECT  1093.28 540.44 1094.3 651.975 ;
     RECT  1094.3 540.44 1094.78 652.36 ;
     RECT  1087.75 662.24 1094.78 1524.28 ;
     RECT  1094.78 540.44 1095.74 1524.28 ;
     RECT  1093.06 1539.2 1095.755 1539.4 ;
     RECT  1085 -70 1098.38 180 ;
     RECT  1095.74 538.76 1098.62 1524.28 ;
     RECT  1098.38 -70 1098.82 181.12 ;
     RECT  1098.62 538.76 1099.525 1526.8 ;
     RECT  1099.525 538.76 1100.06 1456.24 ;
     RECT  1100.06 538.34 1100.26 1456.24 ;
     RECT  1100.26 538.34 1100.74 1376.02 ;
     RECT  1099.525 1466.96 1101.02 1526.8 ;
     RECT  1095.755 1538.61 1101.02 1539.4 ;
     RECT  1093.06 1548.02 1101.5 1549.06 ;
     RECT  1100.74 538.34 1102.46 1065.64 ;
     RECT  1100.26 1384.64 1103.62 1456.24 ;
     RECT  1103.62 1409 1103.7 1456.24 ;
     RECT  1103.7 1409 1104.1 1452.63 ;
     RECT  1101.02 1466.96 1104.1 1539.4 ;
     RECT  1103.62 1384.64 1104.365 1399.54 ;
     RECT  1104.1 1467.345 1105.06 1539.4 ;
     RECT  1104.1 1428.74 1105.12 1452.63 ;
     RECT  1105.06 1467.345 1105.12 1526.8 ;
     RECT  1104.365 1384.64 1105.14 1398.7 ;
     RECT  1105.12 1490.48 1105.14 1515.88 ;
     RECT  1105.06 1539.2 1105.54 1539.4 ;
     RECT  1100.74 1076.78 1106.02 1376.02 ;
     RECT  1104.1 1409 1106.02 1418.86 ;
     RECT  1105.12 1428.74 1106.02 1451.62 ;
     RECT  1105.12 1467.38 1106.02 1481.86 ;
     RECT  1105.14 1490.48 1106.02 1493.62 ;
     RECT  1105.14 1504.34 1106.02 1515.88 ;
     RECT  1106.02 1490.48 1106.5 1490.68 ;
     RECT  1101.5 223.76 1107.46 223.96 ;
     RECT  1105.14 1384.64 1107.46 1394.5 ;
     RECT  1101.5 1548.02 1107.46 1554.94 ;
     RECT  1102.46 532.88 1109.18 1065.64 ;
     RECT  1109.18 531.62 1110.08 1065.64 ;
     RECT  1107.46 1384.64 1110.62 1388.62 ;
     RECT  1106.02 1076.78 1112.06 1371.4 ;
     RECT  1112.06 1075.94 1112.26 1371.4 ;
     RECT  1105.12 1526.6 1112.74 1526.8 ;
     RECT  1112.26 1108.28 1114.46 1371.4 ;
     RECT  1110.62 1382.54 1114.46 1388.62 ;
     RECT  1107.46 1554.74 1115.14 1554.94 ;
     RECT  1112.26 1075.94 1115.18 1094.79 ;
     RECT  1110.08 530.61 1115.9 1065.64 ;
     RECT  1115.18 1075.1 1115.9 1094.79 ;
     RECT  1114.46 1108.28 1115.9 1388.62 ;
     RECT  1082.5 1582.04 1116.58 1582.24 ;
     RECT  1116.38 1414.46 1117.06 1414.66 ;
     RECT  1115.9 530.61 1117.735 1094.79 ;
     RECT  1115.9 1108.28 1120.16 1389.04 ;
     RECT  1117.735 526.58 1121.18 1094.79 ;
     RECT  1120.16 1108.28 1121.18 1389.63 ;
     RECT  1121.18 526.58 1122.62 1095.46 ;
     RECT  1121.18 1108.28 1122.62 1391.98 ;
     RECT  1122.62 526.58 1125.98 1391.98 ;
     RECT  1125.98 526.58 1127.19 1393.24 ;
     RECT  1127.19 215.36 1132.81 1583.92 ;
     RECT  1132.81 519.02 1139.62 1388.62 ;
     RECT  1098.82 -70 1139.9 180 ;
     RECT  1085 1620 1139.9 1870 ;
     RECT  1139.9 -70 1140.1 181.12 ;
     RECT  1139.62 519.86 1140.1 1388.62 ;
     RECT  1139.9 1619.42 1140.1 1870 ;
     RECT  1140.1 519.86 1150.18 1386.1 ;
     RECT  1150.18 519.86 1151.9 1385.26 ;
     RECT  1140.1 -70 1155 180 ;
     RECT  1140.1 1620 1155 1870 ;
     RECT  1151.9 519.02 1155.26 1385.26 ;
     RECT  1155.26 518.6 1159.3 1385.26 ;
     RECT  1155 0 1173 180 ;
     RECT  1155 1620 1173 1800 ;
     RECT  1159.3 518.6 1173.22 1384.84 ;
     RECT  1173.22 519.02 1173.5 1384.84 ;
     RECT  1173.5 519.02 1173.98 1388.62 ;
     RECT  1173.98 519.02 1175.9 1393.24 ;
     RECT  1175.9 519.02 1176.38 1393.66 ;
     RECT  1176.38 519.02 1183.58 1400.8 ;
     RECT  1182.14 223.76 1195.19 223.96 ;
     RECT  1162.46 507.26 1195.19 507.46 ;
     RECT  1183.58 519.02 1195.19 1401.22 ;
     RECT  1195.19 219.14 1200.81 1580.14 ;
     RECT  1200.81 609.32 1202.98 1393.24 ;
     RECT  1202.98 677.36 1204.9 1393.24 ;
     RECT  1204.9 677.36 1205.38 1373.71 ;
     RECT  1205.38 1373.51 1205.62 1373.71 ;
     RECT  1200.81 534.14 1209.98 600.28 ;
     RECT  1202.98 609.32 1209.98 668.74 ;
     RECT  1173 1620 1209.98 1870 ;
     RECT  1205.38 677.36 1211.14 1364.26 ;
     RECT  1209.98 534.14 1212.38 668.74 ;
     RECT  1211.14 677.36 1212.38 1363.42 ;
     RECT  1212.38 534.14 1214.5 1363.42 ;
     RECT  1214.5 644.01 1216.42 1363.42 ;
     RECT  1214.5 534.14 1218.34 633.46 ;
     RECT  1216.42 1311.56 1223.14 1363.42 ;
     RECT  1223.14 1311.56 1223.62 1361.74 ;
     RECT  1200.81 507.26 1223.9 507.46 ;
     RECT  1204.9 1388.42 1223.9 1393.24 ;
     RECT  1223.9 506.84 1224.1 507.46 ;
     RECT  1216.42 644.01 1224.58 1302.94 ;
     RECT  1218.34 542.12 1226.78 633.46 ;
     RECT  1224.58 644.01 1226.78 1302.53 ;
     RECT  1223.9 1386.32 1228.42 1393.24 ;
     RECT  1223.62 1313.24 1231.3 1361.74 ;
     RECT  1226.78 542.12 1233.605 1302.53 ;
     RECT  1231.3 1317.02 1234.18 1361.74 ;
     RECT  1233.605 542.12 1236.1 1301.68 ;
     RECT  1236.1 542.12 1237.54 1294.96 ;
     RECT  1234.18 1320.38 1237.54 1361.74 ;
     RECT  1237.54 542.12 1238.5 542.32 ;
     RECT  1237.54 1346.42 1238.5 1361.74 ;
     RECT  1237.54 1320.38 1239.46 1337.38 ;
     RECT  1237.54 556.82 1240.42 1294.96 ;
     RECT  1240.42 557.24 1240.9 1294.96 ;
     RECT  1240.9 557.625 1241.38 1294.96 ;
     RECT  1241.38 557.625 1241.41 1289.92 ;
     RECT  1241.41 557.66 1241.86 1289.92 ;
     RECT  1173 -70 1243 180 ;
     RECT  1209.98 1616.06 1243 1870 ;
     RECT  1241.86 557.66 1244.74 1288.66 ;
     RECT  1248.38 534.98 1249.28 536.02 ;
     RECT  1224.1 506.84 1249.34 507.04 ;
     RECT  1248.86 456.02 1249.76 456.22 ;
     RECT  1248.86 471.14 1249.76 473.44 ;
     RECT  1249.28 534.945 1249.82 536.02 ;
     RECT  1249.34 506.84 1250.24 511.66 ;
     RECT  1249.82 531.62 1250.72 539.38 ;
     RECT  1249.76 455.01 1250.78 456.22 ;
     RECT  1243.1 496.76 1250.78 497.38 ;
     RECT  1250.78 455.01 1251.26 458.74 ;
     RECT  1249.76 470.13 1251.26 473.44 ;
     RECT  1250.78 486.26 1251.68 497.38 ;
     RECT  1250.24 506.84 1251.74 512.67 ;
     RECT  1251.74 506.84 1252.64 515.86 ;
     RECT  1244.74 557.66 1252.7 1282.36 ;
     RECT  1252.64 506.84 1253.18 515.895 ;
     RECT  1250.72 530.61 1253.18 539.38 ;
     RECT  1252.7 554.3 1253.6 1282.36 ;
     RECT  1253.18 506.84 1253.66 516.28 ;
     RECT  1251.26 455.01 1254.14 473.44 ;
     RECT  1254.14 455.01 1254.62 474.28 ;
     RECT  1251.68 485.25 1254.62 497.38 ;
     RECT  1253.66 506.84 1254.62 517.12 ;
     RECT  1253.18 526.58 1254.62 539.38 ;
     RECT  1253.6 553.29 1254.62 1282.36 ;
     RECT  1254.62 526.58 1255.78 1287.82 ;
     RECT  1254.62 455.01 1255.95 517.12 ;
     RECT  1255.95 451.4 1256.06 517.12 ;
     RECT  1255.78 526.58 1256.06 600.28 ;
     RECT  1255.78 609.32 1256.49 1287.82 ;
     RECT  1256.06 451.4 1256.54 600.28 ;
     RECT  1256.49 1079.72 1257.5 1287.82 ;
     RECT  1256.49 609.32 1257.7 1069 ;
     RECT  1258.46 1302.74 1259.36 1302.94 ;
     RECT  1257.5 1079.72 1259.9 1291.18 ;
     RECT  1243 0 1261 180 ;
     RECT  1243 1616.06 1261 1800 ;
     RECT  1259.9 1079.72 1261.06 1292.86 ;
     RECT  1261.06 1080.56 1261.82 1292.86 ;
     RECT  1259.36 1301.73 1261.82 1302.94 ;
     RECT  1261.82 1080.56 1263.26 1302.94 ;
     RECT  1263.26 1080.56 1264.16 1305.46 ;
     RECT  1257.7 609.32 1264.9 1068.16 ;
     RECT  1264.9 1015.04 1265.38 1068.16 ;
     RECT  1265.38 1015.04 1266.325 1067.74 ;
     RECT  1264.16 1080.56 1266.34 1306.47 ;
     RECT  1266.34 1099.04 1266.62 1306.47 ;
     RECT  1256.54 450.98 1267.1 600.28 ;
     RECT  1264.9 609.32 1267.1 1006.42 ;
     RECT  1267.1 450.98 1269.02 1006.42 ;
     RECT  1266.325 1015.04 1269.7 1066.9 ;
     RECT  1269.7 1015.04 1270.18 1063.96 ;
     RECT  1270.18 1015.04 1270.66 1031.2 ;
     RECT  1270.18 1040.24 1270.66 1063.96 ;
     RECT  1270.46 222.08 1270.94 222.28 ;
     RECT  1270.66 1040.24 1271.62 1043.38 ;
     RECT  1266.62 1099.04 1272.38 1313.44 ;
     RECT  1266.34 1080.56 1273.06 1088.32 ;
     RECT  1269.02 446.78 1273.82 1006.42 ;
     RECT  1270.66 1015.04 1273.82 1030.37 ;
     RECT  1261 1616.06 1274.5 1870 ;
     RECT  1273.06 1085.6 1275.26 1088.32 ;
     RECT  1272.38 1099.04 1275.26 1313.86 ;
     RECT  1270.94 222.08 1276.42 223.96 ;
     RECT  1261 -70 1277.42 180 ;
     RECT  1277.42 -70 1277.86 180.7 ;
     RECT  1276.42 223.76 1277.86 223.96 ;
     RECT  1238.5 1354.4 1277.86 1361.74 ;
     RECT  1273.82 446.78 1279.685 1030.37 ;
     RECT  1279.685 446.78 1281.02 1030.36 ;
     RECT  1275.26 1085.6 1281.98 1313.86 ;
     RECT  1281.02 440.48 1282.18 1030.36 ;
     RECT  1282.18 440.48 1282.94 1027.84 ;
     RECT  1281.98 1083.5 1282.94 1313.86 ;
     RECT  1271.62 1043.18 1284.38 1043.38 ;
     RECT  1270.66 1052.84 1284.38 1063.96 ;
     RECT  1282.94 439.64 1285.28 1027.84 ;
     RECT  1285.28 436.665 1286.3 1027.84 ;
     RECT  1284.38 1043.18 1286.5 1063.96 ;
     RECT  1286.5 1043.18 1286.78 1062.7 ;
     RECT  1282.94 1080.14 1286.78 1313.86 ;
     RECT  1239.46 1322.48 1286.78 1337.38 ;
     RECT  1286.78 1078.04 1288.9 1337.38 ;
     RECT  1286.3 436.28 1289.86 1027.84 ;
     RECT  1286.78 1041.5 1290.34 1062.7 ;
     RECT  1289.86 436.28 1293.98 658.66 ;
     RECT  1290.34 1041.5 1296.38 1045.06 ;
     RECT  1296.38 1038.56 1297.34 1045.06 ;
     RECT  1297.34 1038.14 1298.24 1045.06 ;
     RECT  1293.98 432.5 1298.78 658.66 ;
     RECT  1289.86 668.12 1298.78 1027.84 ;
     RECT  1298.24 1037.13 1301.18 1045.06 ;
     RECT  1301.18 1037.13 1301.38 1045.48 ;
     RECT  1301.38 1037.13 1303.3 1044.64 ;
     RECT  1288.9 1078.04 1303.58 1317.64 ;
     RECT  1288.9 1326.26 1303.58 1337.38 ;
     RECT  1298.78 432.5 1304 1027.84 ;
     RECT  1304 432.33 1306.94 1027.84 ;
     RECT  1306.94 432.33 1309.06 1028.26 ;
     RECT  1309.06 679.46 1309.34 1028.26 ;
     RECT  1303.3 1037.13 1309.34 1043.38 ;
     RECT  1309.06 432.33 1311.445 667.48 ;
     RECT  1309.34 679.46 1312.185 1043.38 ;
     RECT  1303.58 1078.04 1312.22 1337.38 ;
     RECT  1228.42 1386.32 1316.26 1392.82 ;
     RECT  1312.185 679.46 1317.5 1045.06 ;
     RECT  1311.445 432.92 1318.18 667.48 ;
     RECT  1318.18 433.34 1318.94 667.48 ;
     RECT  1317.5 678.2 1318.94 1045.06 ;
     RECT  1312.22 1075.1 1319.36 1337.38 ;
     RECT  1318.94 433.34 1320.1 1045.06 ;
     RECT  1320.1 437.54 1321.1 1045.06 ;
     RECT  1321.1 437.54 1321.34 1045.9 ;
     RECT  1290.34 1054.94 1321.34 1062.7 ;
     RECT  1319.36 1074.93 1323.26 1337.38 ;
     RECT  1323.26 1071.74 1324.16 1337.38 ;
     RECT  1321.34 437.54 1329.02 1062.7 ;
     RECT  1329.02 433.76 1329.5 1062.7 ;
     RECT  1329.5 432.92 1330.46 1062.7 ;
     RECT  1324.16 1071.705 1330.46 1337.38 ;
     RECT  1277.86 -70 1331 180 ;
     RECT  1274.5 1620 1331 1870 ;
     RECT  1330.46 432.92 1331.19 1337.38 ;
     RECT  1277.86 1354.4 1331.19 1356.7 ;
     RECT  1316.26 1386.32 1331.19 1386.52 ;
     RECT  1331.19 215.36 1336.81 1583.92 ;
     RECT  1336.81 432.5 1338.82 1337.38 ;
     RECT  1338.82 432.92 1339.3 1337.38 ;
     RECT  1331 0 1349 180 ;
     RECT  1331 1620 1349 1800 ;
     RECT  1339.3 433.34 1351.1 1337.38 ;
     RECT  1351.1 432.92 1352.74 1337.38 ;
     RECT  1352.74 432.92 1353.5 732.58 ;
     RECT  1352.74 742.29 1353.685 1337.38 ;
     RECT  1353.5 432.08 1355.14 732.58 ;
     RECT  1355.14 432.92 1358.02 732.58 ;
     RECT  1353.685 742.46 1358.02 1337.38 ;
     RECT  1358.3 222.08 1358.78 222.28 ;
     RECT  1336.81 1354.4 1359.26 1356.7 ;
     RECT  1358.02 948.26 1360.42 1337.38 ;
     RECT  1349 -70 1362.38 180 ;
     RECT  1358.78 222.08 1364.26 223.96 ;
     RECT  1358.02 742.46 1365.02 937.96 ;
     RECT  1365.02 741.62 1365.22 937.96 ;
     RECT  1358.02 435.86 1365.5 732.58 ;
     RECT  1365.22 741.62 1365.5 901.42 ;
     RECT  1364.26 223.76 1365.7 223.96 ;
     RECT  1359.26 1354.4 1365.7 1363.42 ;
     RECT  1362.38 -70 1367.14 180.7 ;
     RECT  1365.22 913.82 1367.42 937.96 ;
     RECT  1365.5 435.86 1368.565 901.42 ;
     RECT  1368.565 826.04 1368.58 901.42 ;
     RECT  1367.42 913.82 1368.86 940.06 ;
     RECT  1360.42 950.36 1368.86 1337.38 ;
     RECT  1368.58 848.13 1369.525 901.42 ;
     RECT  1368.565 435.86 1371.94 817.42 ;
     RECT  1369.525 849.14 1372.9 901.42 ;
     RECT  1372.9 849.56 1373.66 901.42 ;
     RECT  1371.94 786.98 1373.86 814.06 ;
     RECT  1373.66 849.56 1374.505 901.84 ;
     RECT  1373.86 813.86 1374.82 814.06 ;
     RECT  1368.58 827.3 1375.3 838.42 ;
     RECT  1374.505 849.56 1375.58 902.26 ;
     RECT  1368.86 913.82 1375.58 1337.38 ;
     RECT  1375.3 828.56 1376.74 838.42 ;
     RECT  1376.74 832.76 1377.7 834.64 ;
     RECT  1377.7 833.6 1378.66 834.64 ;
     RECT  1371.94 435.86 1381.58 776.68 ;
     RECT  1373.86 786.98 1381.58 803.57 ;
     RECT  1381.58 435.86 1381.82 803.57 ;
     RECT  1381.82 425.78 1382.3 803.57 ;
     RECT  1382.3 425.78 1382.72 803.98 ;
     RECT  1382.72 424.77 1384.22 803.98 ;
     RECT  1384.22 420.74 1388.06 803.98 ;
     RECT  1388.06 420.74 1391.9 811.54 ;
     RECT  1391.9 413.6 1395.74 811.54 ;
     RECT  1375.58 849.56 1396.7 1337.38 ;
     RECT  1395.74 413.6 1399.19 814.06 ;
     RECT  1389.5 827.72 1399.19 827.92 ;
     RECT  1396.7 842 1399.19 1337.38 ;
     RECT  1365.7 1354.4 1399.19 1356.7 ;
     RECT  1336.81 1386.32 1399.19 1386.52 ;
     RECT  1367.14 -70 1403.9 180 ;
     RECT  1349 1620 1403.9 1870 ;
     RECT  1403.9 -70 1404.1 180.7 ;
     RECT  1399.19 219.14 1404.81 1580.14 ;
     RECT  1404.81 1386.32 1405.54 1386.52 ;
     RECT  1403.9 1619.42 1405.54 1870 ;
     RECT  1404.81 827.72 1406.02 827.92 ;
     RECT  1404.81 855.02 1406.5 856.9 ;
     RECT  1406.5 855.44 1409.86 856.9 ;
     RECT  1404.81 867.2 1413.53 1337.38 ;
     RECT  1404.81 413.18 1414.66 810.7 ;
     RECT  1404.81 842 1414.855 842.2 ;
     RECT  1414.855 841.16 1414.94 842.2 ;
     RECT  1414.94 840.32 1415.815 842.2 ;
     RECT  1415.815 833.6 1415.9 842.2 ;
     RECT  1415.9 832.76 1416.295 842.2 ;
     RECT  1414.66 414.02 1418.005 810.7 ;
     RECT  1409.86 855.44 1418.78 855.64 ;
     RECT  1413.53 866.86 1418.78 1337.38 ;
     RECT  1404.1 -70 1419 180 ;
     RECT  1405.54 1620 1419 1870 ;
     RECT  1416.295 829.4 1421.095 842.2 ;
     RECT  1418.005 416.54 1421.18 810.7 ;
     RECT  1421.095 821.84 1421.18 842.2 ;
     RECT  1418.78 855.44 1422.535 1337.38 ;
     RECT  1421.18 416.54 1422.82 842.2 ;
     RECT  1422.82 416.54 1425.22 489.4 ;
     RECT  1422.82 498.02 1426.94 842.2 ;
     RECT  1422.535 851.66 1426.94 1337.38 ;
     RECT  1425.22 417.21 1427.14 489.4 ;
     RECT  1426.94 498.02 1431.74 1337.38 ;
     RECT  1427.14 417.21 1433.66 487.3 ;
     RECT  1433.66 413.18 1436.06 487.3 ;
     RECT  1431.74 496.34 1436.06 1337.38 ;
     RECT  1419 0 1437 180 ;
     RECT  1419 1620 1437 1800 ;
     RECT  1436.06 413.18 1437.22 1337.38 ;
     RECT  1437.22 413.6 1444.9 1337.38 ;
     RECT  1444.9 417.21 1447.765 1337.38 ;
     RECT  1447.765 802.1 1448.26 1337.38 ;
     RECT  1447.765 417.21 1449.155 792.655 ;
     RECT  1449.155 417.21 1449.22 791.82 ;
     RECT  1449.22 787.385 1449.605 791.82 ;
     RECT  1448.26 802.1 1450.66 811.12 ;
     RECT  1448.26 821 1450.66 1337.38 ;
     RECT  1449.22 417.21 1451.14 778.36 ;
     RECT  1450.66 802.1 1451.14 806.08 ;
     RECT  1451.14 417.21 1452.1 777.94 ;
     RECT  1450.66 822.26 1452.1 1337.38 ;
     RECT  1452.1 824.36 1453.54 1337.38 ;
     RECT  1453.54 824.78 1454.5 1337.38 ;
     RECT  1454.5 824.78 1455.7 860.68 ;
     RECT  1452.1 417.21 1455.925 777.27 ;
     RECT  1455.7 828.56 1455.94 860.68 ;
     RECT  1455.925 417.21 1456.7 775.84 ;
     RECT  1455.94 851.66 1456.9 860.68 ;
     RECT  1456.9 851.66 1457.38 851.86 ;
     RECT  1454.5 871.4 1457.38 1337.38 ;
     RECT  1455.94 828.56 1457.86 841.36 ;
     RECT  1456.7 413.6 1459.3 775.84 ;
     RECT  1457.86 828.56 1459.3 834.64 ;
     RECT  1457.38 874.34 1462.66 1337.38 ;
     RECT  1449.605 787.385 1463.555 789.28 ;
     RECT  1463.555 788.22 1464.005 789.28 ;
     RECT  1464.005 788.24 1464.58 789.28 ;
     RECT  1462.66 878.96 1464.58 1337.38 ;
     RECT  1459.3 413.6 1464.81 773.32 ;
     RECT  1464.81 770.18 1466.98 773.32 ;
     RECT  1464.58 883.58 1467.46 1337.38 ;
     RECT  1467.46 889.04 1467.94 896.8 ;
     RECT  1464.81 413.6 1468.42 761.56 ;
     RECT  1467.94 889.46 1468.42 893.44 ;
     RECT  1451.14 802.1 1468.9 802.3 ;
     RECT  1468.42 893.24 1468.9 893.44 ;
     RECT  1468.42 413.6 1471.58 758.62 ;
     RECT  1471.58 413.18 1472.26 758.62 ;
     RECT  1467.46 911.72 1472.74 1337.38 ;
     RECT  1472.74 912.56 1473.22 1337.38 ;
     RECT  1472.26 413.18 1476.58 756.52 ;
     RECT  1473.22 914.66 1478.02 1337.38 ;
     RECT  1476.58 414.02 1479.925 756.52 ;
     RECT  1478.02 914.66 1481.38 1000.54 ;
     RECT  1481.38 915.92 1481.86 1000.54 ;
     RECT  1481.86 915.92 1482.34 1000.12 ;
     RECT  1482.34 921.38 1483.3 1000.12 ;
     RECT  1478.02 1010.84 1484.97 1056.82 ;
     RECT  1483.3 921.38 1485.185 996.34 ;
     RECT  1485.185 921.38 1486.18 995.08 ;
     RECT  1484.97 1010.84 1486.46 1055.56 ;
     RECT  1468.7 775.22 1486.66 775.42 ;
     RECT  1486.46 1009.16 1489.06 1055.56 ;
     RECT  1489.06 1009.16 1490.5 1051.78 ;
     RECT  1478.02 1066.7 1491.94 1337.38 ;
     RECT  1486.18 921.38 1492.185 994.66 ;
     RECT  1490.5 1010.42 1492.42 1051.78 ;
     RECT  1492.42 1010.42 1492.9 1049.26 ;
     RECT  1492.9 1019.66 1494.34 1048.84 ;
     RECT  1479.925 418.64 1494.62 756.52 ;
     RECT  1494.34 1019.66 1495.3 1031.2 ;
     RECT  1495.3 1019.66 1495.78 1030.36 ;
     RECT  1494.34 1042.34 1495.78 1048.84 ;
     RECT  1495.78 1025.96 1496.26 1030.36 ;
     RECT  1495.78 1044.86 1496.26 1048.84 ;
     RECT  1496.26 1028.48 1496.74 1030.36 ;
     RECT  1464.58 788.24 1497.02 788.44 ;
     RECT  1496.74 1028.9 1497.22 1030.36 ;
     RECT  1492.185 920.54 1497.5 994.66 ;
     RECT  1497.22 1028.9 1497.7 1029.1 ;
     RECT  1496.26 1045.7 1497.7 1048.84 ;
     RECT  1494.62 418.22 1498.825 756.52 ;
     RECT  1491.94 1067.12 1499.14 1337.38 ;
     RECT  1498.825 418.22 1499.32 757.375 ;
     RECT  1499.32 418.22 1501.28 758.21 ;
     RECT  1497.02 781.1 1501.54 788.44 ;
     RECT  1501.28 417.21 1503.26 758.21 ;
     RECT  1501.54 788.24 1504.42 788.44 ;
     RECT  1497.5 920.54 1504.9 996.34 ;
     RECT  1504.9 928.52 1505.38 996.34 ;
     RECT  1505.38 930.2 1505.86 996.34 ;
     RECT  1505.86 931.88 1505.95 996.34 ;
     RECT  1505.95 931.88 1505.955 996.13 ;
     RECT  1505.955 931.88 1506.6 995.92 ;
     RECT  1506.6 931.88 1506.82 995.08 ;
     RECT  1437 -70 1507 180 ;
     RECT  1437 1620 1507 1870 ;
     RECT  1503.26 417.21 1507.3 758.62 ;
     RECT  1506.82 931.88 1507.3 994.66 ;
     RECT  1499.14 1067.54 1507.78 1337.38 ;
     RECT  1507.3 417.21 1508.725 756.52 ;
     RECT  1507.3 939.44 1510.66 994.66 ;
     RECT  1508.725 417.38 1511.14 756.52 ;
     RECT  1511.14 417.38 1512.1 753.58 ;
     RECT  1510.66 951.62 1512.1 994.66 ;
     RECT  1507.78 1071.74 1512.1 1337.38 ;
     RECT  1512.1 951.62 1512.34 951.82 ;
     RECT  1512.1 1075.94 1512.58 1337.38 ;
     RECT  1512.58 1075.94 1513.06 1108.06 ;
     RECT  1512.1 421.16 1514.02 753.58 ;
     RECT  1512.1 962.12 1514.5 994.66 ;
     RECT  1512.58 1117.1 1514.98 1337.38 ;
     RECT  1514.5 962.12 1515.94 989.2 ;
     RECT  1513.06 1075.94 1516.42 1106.38 ;
     RECT  1515.94 964.64 1517.38 989.2 ;
     RECT  1514.98 1117.1 1517.86 1137.04 ;
     RECT  1517.86 1128.42 1518.245 1137.04 ;
     RECT  1517.38 964.64 1518.82 988.36 ;
     RECT  1516.42 1075.94 1519.285 1105.54 ;
     RECT  1519.285 1075.94 1519.3 1100.5 ;
     RECT  1518.82 964.64 1519.78 982.9 ;
     RECT  1519.3 1075.94 1520.74 1076.14 ;
     RECT  1517.86 1117.1 1522.18 1118.14 ;
     RECT  1518.245 1128.44 1522.18 1137.04 ;
     RECT  1519.78 979.76 1522.66 982.9 ;
     RECT  1519.3 1089.38 1522.66 1100.5 ;
     RECT  1522.66 979.76 1523.14 980.8 ;
     RECT  1514.02 421.16 1523.9 751.9 ;
     RECT  1522.66 1089.38 1524.58 1090.84 ;
     RECT  1523.9 418.22 1524.8 751.9 ;
     RECT  1507 0 1525 180 ;
     RECT  1507 1620 1525 1800 ;
     RECT  1522.18 1128.44 1526.02 1133.26 ;
     RECT  1404.81 1354.4 1526.3 1356.7 ;
     RECT  1524.8 417.21 1528.22 751.9 ;
     RECT  1528.22 416.54 1529.66 751.9 ;
     RECT  1529.66 416.54 1530.62 754 ;
     RECT  1526.02 1133.06 1531.58 1133.26 ;
     RECT  1530.62 416.54 1533.02 754.84 ;
     RECT  1533.02 414.02 1535.19 754.84 ;
     RECT  1459.3 834.44 1535.19 834.64 ;
     RECT  1529.66 889.04 1535.19 889.24 ;
     RECT  1519.78 964.64 1535.19 964.84 ;
     RECT  1534.46 1058.3 1535.19 1058.5 ;
     RECT  1522.66 1099.46 1535.19 1100.5 ;
     RECT  1522.94 1115.84 1535.19 1116.04 ;
     RECT  1531.58 1133.06 1535.19 1137.46 ;
     RECT  1514.98 1146.08 1535.19 1337.38 ;
     RECT  1526.3 1354.4 1535.19 1360.9 ;
     RECT  1535.19 215.36 1540.81 1583.92 ;
     RECT  1540.81 1137.26 1540.9 1147.54 ;
     RECT  1540.81 889.04 1541.38 889.24 ;
     RECT  1540.81 1173.21 1541.38 1221.88 ;
     RECT  1541.38 1173.21 1541.845 1208.19 ;
     RECT  1540.81 1159.1 1541.86 1163.5 ;
     RECT  1541.845 1174.64 1542.325 1208.19 ;
     RECT  1541.38 1220.42 1542.34 1221.88 ;
     RECT  1540.81 1231.34 1542.34 1258 ;
     RECT  1541.86 1163.3 1542.82 1163.5 ;
     RECT  1542.34 1231.34 1542.82 1242.88 ;
     RECT  1542.34 1252.76 1542.82 1258 ;
     RECT  1540.81 1058.3 1543.3 1058.5 ;
     RECT  1542.82 1237.63 1543.3 1242.88 ;
     RECT  1542.82 1252.76 1543.78 1253.38 ;
     RECT  1540.81 1325.84 1544.26 1337.38 ;
     RECT  1542.325 1174.64 1544.74 1208.02 ;
     RECT  1540.81 413.18 1545.22 750.22 ;
     RECT  1544.74 1174.64 1545.22 1192.9 ;
     RECT  1544.74 1202.78 1545.22 1208.02 ;
     RECT  1545.22 1207.4 1545.7 1208.02 ;
     RECT  1543.3 1237.63 1546.085 1239.94 ;
     RECT  1540.81 1099.46 1546.66 1100.5 ;
     RECT  1546.085 1237.64 1546.66 1239.94 ;
     RECT  1545.22 598.82 1547.62 750.22 ;
     RECT  1540.81 1354.4 1547.62 1360.9 ;
     RECT  1540.9 1137.26 1548.1 1144.6 ;
     RECT  1545.22 413.18 1549.06 589.36 ;
     RECT  1547.62 599.24 1550.3 750.22 ;
     RECT  1540.81 1029.32 1551.94 1029.52 ;
     RECT  1550.3 599.24 1552.22 750.64 ;
     RECT  1545.22 1180.505 1552.355 1192.9 ;
     RECT  1552.355 1181.34 1552.805 1192.9 ;
     RECT  1552.805 1186.4 1553.38 1192.9 ;
     RECT  1540.81 1119.62 1555.1 1119.82 ;
     RECT  1548.1 1144.4 1555.3 1144.6 ;
     RECT  1549.06 414.02 1556.54 589.36 ;
     RECT  1552.22 599.24 1556.54 751.06 ;
     RECT  1540.81 863.84 1558.66 864.04 ;
     RECT  1551.74 972.2 1558.66 972.4 ;
     RECT  1556.54 414.02 1559.14 751.06 ;
     RECT  1559.14 418.64 1560.58 751.06 ;
     RECT  1560.58 451.785 1561.06 751.06 ;
     RECT  1561.06 451.785 1561.09 747.03 ;
     RECT  1560.58 418.64 1561.3 440.26 ;
     RECT  1561.3 420.74 1562.5 440.26 ;
     RECT  1561.09 451.82 1562.5 747.03 ;
     RECT  1540.81 1280.9 1565.66 1293.28 ;
     RECT  1558.46 928.94 1565.86 929.14 ;
     RECT  1555.1 1115.84 1565.86 1119.82 ;
     RECT  1565.66 1274.6 1565.86 1293.28 ;
     RECT  1562.5 420.74 1566.275 437.335 ;
     RECT  1566.275 420.74 1566.725 436.5 ;
     RECT  1562.5 451.82 1568.245 713.26 ;
     RECT  1566.725 420.74 1568.26 428.5 ;
     RECT  1540.81 1378.76 1569.5 1378.96 ;
     RECT  1565.86 1293.08 1569.7 1293.28 ;
     RECT  1569.5 1378.76 1569.7 1385.68 ;
     RECT  1562.5 722.72 1571.14 747.03 ;
     RECT  1568.245 455.18 1573.06 713.26 ;
     RECT  1565.66 1065.44 1573.06 1065.64 ;
     RECT  1553.38 1186.4 1573.06 1190.38 ;
     RECT  1573.06 455.18 1573.54 511.66 ;
     RECT  1573.06 523.64 1573.54 713.26 ;
     RECT  1571.14 722.72 1573.54 738.88 ;
     RECT  1551.26 1010.42 1573.82 1010.62 ;
     RECT  1573.54 466.1 1574.5 505.11 ;
     RECT  1546.66 1239.74 1574.5 1239.94 ;
     RECT  1573.54 455.18 1574.98 455.38 ;
     RECT  1574.5 469.88 1574.98 486.04 ;
     RECT  1573.54 722.72 1574.98 735.52 ;
     RECT  1544.26 1325.84 1574.98 1328.56 ;
     RECT  1573.54 527 1575.46 713.26 ;
     RECT  1573.06 1186.4 1575.74 1189.96 ;
     RECT  1574.98 469.88 1575.94 484.78 ;
     RECT  1574.98 722.72 1575.94 722.92 ;
     RECT  1569.5 1264.52 1575.94 1264.72 ;
     RECT  1575.46 527 1576.42 706.54 ;
     RECT  1575.74 1512.74 1576.42 1512.94 ;
     RECT  1558.46 802.52 1576.7 802.72 ;
     RECT  1565.86 1274.6 1576.7 1281.1 ;
     RECT  1547.62 1354.4 1576.7 1356.7 ;
     RECT  1574.5 496.76 1576.9 505.11 ;
     RECT  1576.42 527 1576.9 554.92 ;
     RECT  1576.42 565.22 1576.9 706.54 ;
     RECT  1574.98 734.9 1576.9 735.52 ;
     RECT  1576.7 800.42 1576.9 802.72 ;
     RECT  1574.98 1328.36 1576.9 1328.56 ;
     RECT  1544.26 1337.18 1576.9 1337.38 ;
     RECT  1576.7 1354.4 1576.9 1365.94 ;
     RECT  1576.9 535.82 1577.38 554.92 ;
     RECT  1576.9 527 1577.86 527.2 ;
     RECT  1540.81 834.44 1578.14 834.64 ;
     RECT  1546.66 1100.3 1578.14 1100.5 ;
     RECT  1577.66 998.66 1578.34 998.86 ;
     RECT  1576.7 1259.9 1578.34 1263.46 ;
     RECT  1577.38 538.17 1578.805 554.92 ;
     RECT  1576.9 565.22 1578.82 706.12 ;
     RECT  1578.14 1086.02 1578.82 1086.22 ;
     RECT  1578.14 1339.7 1578.82 1339.9 ;
     RECT  1575.94 474.5 1579.3 484.78 ;
     RECT  1572.86 979.34 1583.9 979.54 ;
     RECT  1575.74 1183.88 1583.9 1189.96 ;
     RECT  1542.34 1220.42 1587.26 1220.62 ;
     RECT  1576.7 397.64 1588.14 397.84 ;
     RECT  1583.9 445.94 1588.14 446.14 ;
     RECT  1579.3 474.5 1588.14 474.7 ;
     RECT  1576.9 497.18 1588.14 505.11 ;
     RECT  1578.805 539.6 1588.14 554.92 ;
     RECT  1578.82 565.22 1588.14 609.52 ;
     RECT  1578.82 620.66 1588.14 706.12 ;
     RECT  1576.9 734.9 1588.14 735.1 ;
     RECT  1574.78 749.6 1588.14 749.8 ;
     RECT  1576.9 800.42 1588.14 800.62 ;
     RECT  1578.14 834.44 1588.14 838 ;
     RECT  1578.62 925.58 1588.14 925.78 ;
     RECT  1583.9 978.5 1588.14 979.54 ;
     RECT  1573.82 1010.42 1588.14 1013.98 ;
     RECT  1587.26 1076.36 1588.14 1076.56 ;
     RECT  1578.14 1100.3 1588.14 1101.76 ;
     RECT  1565.86 1119.62 1588.14 1119.82 ;
     RECT  1583.9 1183.88 1588.14 1197.94 ;
     RECT  1587.26 1220.42 1588.14 1228.18 ;
     RECT  1587.74 1244.36 1588.14 1244.56 ;
     RECT  1578.34 1259.9 1588.14 1260.1 ;
     RECT  1576.7 1274.18 1588.14 1281.1 ;
     RECT  1576.7 1317.86 1588.14 1318.06 ;
     RECT  1576.9 1361.96 1588.14 1365.94 ;
     RECT  1569.7 1385.48 1588.14 1385.68 ;
     RECT  1525 -70 1595 180 ;
     RECT  1525 1620 1595 1870 ;
     RECT  1588.14 215.36 1597.86 1583.92 ;
     RECT  1595 0 1620 180 ;
     RECT  1597.86 219.14 1620 1580.14 ;
     RECT  1595 1620 1620 1800 ;
     RECT  1620 0 1800 1800 ;
     RECT  1800 205 1870 275 ;
     RECT  1800 293 1870 363 ;
     RECT  1800 381 1870 451 ;
     RECT  1800 469 1870 539 ;
     RECT  1800 557 1870 627 ;
     RECT  1800 645 1870 715 ;
     RECT  1800 733 1870 803 ;
     RECT  1800 821 1870 891 ;
     RECT  1800 909 1870 979 ;
     RECT  1800 997 1870 1067 ;
     RECT  1800 1085 1870 1155 ;
     RECT  1800 1173 1870 1243 ;
     RECT  1800 1261 1870 1331 ;
     RECT  1800 1349 1870 1419 ;
     RECT  1800 1437 1870 1507 ;
     RECT  1800 1525 1870 1595 ;
    LAYER Metal3 ;
     RECT  205 -70 275 0 ;
     RECT  293 -70 363 0 ;
     RECT  381 -70 451 0 ;
     RECT  469 -70 539 0 ;
     RECT  557 -70 627 0 ;
     RECT  645 -70 715 0 ;
     RECT  733 -70 803 0 ;
     RECT  821 -70 891 0 ;
     RECT  909 -70 979 0 ;
     RECT  997 -70 1067 0 ;
     RECT  1085 -70 1155 0 ;
     RECT  1173 -70 1243 0 ;
     RECT  1261 -70 1331 0 ;
     RECT  1349 -70 1419 0 ;
     RECT  1437 -70 1507 0 ;
     RECT  1525 -70 1595 0 ;
     RECT  0 0 1800 178 ;
     RECT  0 178 180 180 ;
     RECT  394.225 178 398.02 180 ;
     RECT  435.725 178 438.34 180 ;
     RECT  482.225 178 485.86 180 ;
     RECT  523.725 178 524.26 180 ;
     RECT  570.225 178 573.775 180 ;
     RECT  611.725 178 612.225 180 ;
     RECT  658.225 178 662.02 180 ;
     RECT  699.725 178 700.42 180 ;
     RECT  746.225 178 749.86 180 ;
     RECT  786.62 178 788.225 180 ;
     RECT  834.225 178 837.775 180 ;
     RECT  875.725 178 876.225 180 ;
     RECT  922.225 178 925.775 180 ;
     RECT  963.725 178 964.42 180 ;
     RECT  1010.225 178 1013.86 180 ;
     RECT  1051.725 178 1052.26 180 ;
     RECT  1098.225 178 1101.775 180 ;
     RECT  1139.725 178 1140.225 180 ;
     RECT  1186.225 178 1190.02 180 ;
     RECT  1225.82 178 1228.225 180 ;
     RECT  1274.225 178 1277.86 180 ;
     RECT  1315.725 178 1316.225 180 ;
     RECT  1362.225 178 1367.14 180 ;
     RECT  1403.725 178 1404.225 180 ;
     RECT  1620 178 1800 180 ;
     RECT  1403.9 180 1404.1 180.7 ;
     RECT  482.54 180 485.86 181.96 ;
     RECT  746.54 180 749.86 181.96 ;
     RECT  1189.58 180 1190.02 181.96 ;
     RECT  1012.7 180 1013.86 184.06 ;
     RECT  922.46 180 923.14 187.3 ;
     RECT  438.14 180 438.34 197.92 ;
     RECT  0 180 178 205 ;
     RECT  1622 180 1800 205 ;
     RECT  524.06 180 524.26 215.315 ;
     RECT  922.46 187.3 922.66 215.315 ;
     RECT  834.62 180 837.7 216.2 ;
     RECT  394.46 180 398.02 217.46 ;
     RECT  1013.66 184.06 1013.86 217.46 ;
     RECT  -70 205 178 219.095 ;
     RECT  202.185 215.315 211.815 219.095 ;
     RECT  570.62 180 573.7 219.095 ;
     RECT  786.62 180 786.82 219.095 ;
     RECT  1189.82 181.96 1190.02 219.095 ;
     RECT  1588.185 215.315 1597.815 219.095 ;
     RECT  1622 205 1870 219.095 ;
     RECT  1013.66 217.46 1020.1 220.18 ;
     RECT  658.46 180 662.02 220.82 ;
     RECT  746.78 181.96 749.86 221.24 ;
     RECT  394.46 217.46 403.78 221.44 ;
     RECT  834.62 216.2 843.94 221.44 ;
     RECT  1019.9 220.18 1020.1 221.44 ;
     RECT  746.78 221.24 756.1 221.86 ;
     RECT  1277.66 180 1277.86 222.08 ;
     RECT  1365.5 180 1367.14 222.08 ;
     RECT  482.78 181.96 485.86 223.54 ;
     RECT  922.46 215.315 928.765 223.96 ;
     RECT  1101.5 180 1101.7 223.96 ;
     RECT  1189.82 219.095 1200.765 223.96 ;
     RECT  1270.46 222.08 1277.86 223.96 ;
     RECT  570.62 219.095 588.765 224.38 ;
     RECT  658.46 220.82 668.26 224.8 ;
     RECT  1270.46 223.96 1270.66 224.8 ;
     RECT  1358.3 222.08 1367.14 224.8 ;
     RECT  1052.06 180 1052.26 230.68 ;
     RECT  515.235 215.315 524.26 255.46 ;
     RECT  875.9 180 876.1 263.02 ;
     RECT  570.62 224.38 570.82 270.16 ;
     RECT  -70 219.095 211.815 275 ;
     RECT  1588.185 219.095 1870 275 ;
     RECT  786.62 219.095 792.765 284.44 ;
     RECT  0 275 211.815 293 ;
     RECT  1588.185 275 1800 293 ;
     RECT  405.02 222.08 405.22 327.7 ;
     RECT  658.46 224.8 658.66 334.84 ;
     RECT  482.78 223.54 482.98 341.98 ;
     RECT  394.46 221.44 394.66 349.12 ;
     RECT  611.9 180 612.1 356.26 ;
     RECT  -70 293 211.815 363 ;
     RECT  1588.185 293 1870 363 ;
     RECT  834.62 221.44 834.82 363.82 ;
     RECT  746.78 221.86 746.98 370.96 ;
     RECT  0 363 211.815 381 ;
     RECT  1588.185 363 1800 381 ;
     RECT  875.9 382.94 876.1 384.62 ;
     RECT  904.7 385.88 904.9 386.3 ;
     RECT  297.5 386.72 297.7 387.14 ;
     RECT  964.22 180 964.42 387.56 ;
     RECT  235.58 383.36 235.78 387.98 ;
     RECT  -70 381 211.815 388.4 ;
     RECT  991.235 219.095 996.765 388.4 ;
     RECT  353.66 384.2 353.86 388.82 ;
     RECT  583.235 224.38 588.765 389.24 ;
     RECT  787.235 284.44 792.765 390.5 ;
     RECT  787.235 390.5 794.5 390.92 ;
     RECT  809.18 391.34 809.38 392.18 ;
     RECT  844.7 381.26 844.9 392.18 ;
     RECT  379.235 219.095 384.765 392.6 ;
     RECT  572.54 388.4 572.74 392.6 ;
     RECT  583.235 389.24 594.82 392.6 ;
     RECT  379.235 392.6 387.46 393.02 ;
     RECT  353.66 388.82 357.22 393.44 ;
     RECT  560.06 389.24 560.26 393.44 ;
     RECT  840.86 392.18 844.9 393.44 ;
     RECT  328.22 385.04 328.42 393.86 ;
     RECT  345.5 393.44 357.22 393.86 ;
     RECT  379.235 393.02 390.82 393.86 ;
     RECT  875.9 384.62 884.74 393.86 ;
     RECT  311.235 215.315 316.765 394.28 ;
     RECT  328.22 393.86 357.22 394.28 ;
     RECT  369.98 393.86 390.82 394.28 ;
     RECT  765.98 393.44 766.18 394.28 ;
     RECT  560.06 393.44 561.22 394.48 ;
     RECT  765.98 394.28 767.14 394.48 ;
     RECT  311.235 394.28 357.22 394.7 ;
     RECT  572.54 392.6 594.82 394.7 ;
     RECT  875.9 393.86 888.1 394.7 ;
     RECT  741.5 394.7 742.18 394.9 ;
     RECT  291.74 387.14 297.7 395.12 ;
     RECT  310.46 394.7 357.22 395.12 ;
     RECT  565.34 394.7 594.82 395.12 ;
     RECT  565.34 395.12 595.78 395.32 ;
     RECT  515.235 255.46 520.765 395.54 ;
     RECT  871.1 394.7 888.1 395.54 ;
     RECT  955.1 387.56 964.42 395.54 ;
     RECT  719.235 215.315 724.765 395.96 ;
     RECT  549.98 380.84 550.18 396.8 ;
     RECT  486.62 392.18 486.82 397.22 ;
     RECT  535.1 383.78 535.3 398.48 ;
     RECT  515.235 395.54 522.34 398.9 ;
     RECT  535.1 398.48 539.14 398.9 ;
     RECT  515.235 398.9 539.14 399.74 ;
     RECT  787.235 390.92 798.34 399.74 ;
     RECT  437.18 399.74 437.38 400.16 ;
     RECT  447.26 390.08 447.46 400.16 ;
     RECT  719.235 395.96 730.66 400.16 ;
     RECT  786.62 399.74 798.34 400.16 ;
     RECT  549.98 396.8 553.54 400.36 ;
     RECT  411.26 391.76 411.46 401 ;
     RECT  514.46 399.74 539.14 401.42 ;
     RECT  549.98 400.36 550.18 401.42 ;
     RECT  682.46 401.84 682.66 402.26 ;
     RECT  923.235 223.96 928.765 402.26 ;
     RECT  273.5 395.54 273.7 402.68 ;
     RECT  682.46 402.26 686.02 402.68 ;
     RECT  700.22 180 700.42 402.68 ;
     RECT  780.86 400.16 798.34 403.52 ;
     RECT  809.18 392.18 815.14 403.52 ;
     RECT  411.26 401 421.06 404.36 ;
     RECT  682.46 402.68 700.42 404.36 ;
     RECT  713.66 400.16 730.66 404.36 ;
     RECT  682.46 404.36 730.66 404.98 ;
     RECT  499.58 405.2 499.78 405.62 ;
     RECT  514.46 401.42 550.18 405.62 ;
     RECT  499.58 405.62 550.18 406.04 ;
     RECT  713.66 404.98 730.66 406.88 ;
     RECT  741.98 394.9 742.18 406.88 ;
     RECT  904.7 386.3 910.66 407.3 ;
     RECT  758.78 397.64 764.26 407.72 ;
     RECT  465.5 389.66 465.7 408.14 ;
     RECT  437.18 400.16 447.46 408.56 ;
     RECT  291.74 395.12 357.22 408.98 ;
     RECT  921.98 402.26 928.765 408.98 ;
     RECT  645.98 408.98 646.18 409.4 ;
     RECT  921.98 408.98 938.5 409.4 ;
     RECT  949.82 395.54 964.42 409.4 ;
     RECT  273.5 402.68 275.14 409.82 ;
     RECT  572.54 395.32 594.82 409.82 ;
     RECT  263.9 409.82 275.14 410.24 ;
     RECT  840.86 393.44 849.22 410.66 ;
     RECT  255.74 410.24 275.14 411.08 ;
     RECT  285.02 408.98 357.22 411.08 ;
     RECT  645.98 409.4 648.1 412.76 ;
     RECT  713.66 406.88 742.18 412.76 ;
     RECT  753.02 407.72 764.26 412.76 ;
     RECT  837.98 410.66 849.22 412.76 ;
     RECT  566.78 409.82 594.82 413.18 ;
     RECT  828.38 412.76 849.22 413.18 ;
     RECT  1535.235 215.315 1540.765 413.18 ;
     RECT  460.7 408.14 465.7 413.6 ;
     RECT  477.02 397.22 486.82 413.6 ;
     RECT  498.62 406.04 550.18 413.6 ;
     RECT  609.5 412.76 609.7 413.6 ;
     RECT  780.86 403.52 815.14 413.6 ;
     RECT  825.98 413.18 849.22 413.6 ;
     RECT  1399.235 219.095 1404.765 413.6 ;
     RECT  1414.46 413.18 1414.66 413.6 ;
     RECT  1476.38 413.18 1476.58 413.6 ;
     RECT  368.54 394.28 390.82 414.02 ;
     RECT  404.06 404.36 421.06 414.02 ;
     RECT  780.86 413.6 849.22 414.02 ;
     RECT  865.82 395.54 888.1 414.02 ;
     RECT  1433.66 413.18 1433.86 414.02 ;
     RECT  1444.7 413.6 1444.9 414.02 ;
     RECT  1456.7 413.6 1456.9 414.02 ;
     RECT  1468.22 413.6 1476.58 414.02 ;
     RECT  1535.235 413.18 1548.58 414.02 ;
     RECT  255.74 411.08 357.22 414.44 ;
     RECT  368.54 414.02 421.06 414.44 ;
     RECT  682.46 404.98 702.82 414.86 ;
     RECT  780.86 414.02 888.1 414.86 ;
     RECT  898.94 407.3 910.66 414.86 ;
     RECT  1391.9 413.6 1414.66 414.86 ;
     RECT  1456.7 414.02 1476.58 414.86 ;
     RECT  921.98 409.4 964.42 415.28 ;
     RECT  609.5 413.6 611.62 415.7 ;
     RECT  645.98 412.76 656.74 415.7 ;
     RECT  566.78 413.18 595.78 415.945 ;
     RECT  991.235 388.4 1005.22 415.945 ;
     RECT  645.98 415.7 658.18 416.54 ;
     RECT  669.02 401 669.22 416.54 ;
     RECT  1533.02 414.02 1559.14 416.54 ;
     RECT  235.58 387.98 241.54 416.96 ;
     RECT  255.74 414.44 421.06 416.96 ;
     RECT  645.98 416.54 669.22 416.96 ;
     RECT  680.06 414.86 702.82 416.96 ;
     RECT  645.98 416.96 702.82 417.38 ;
     RECT  713.66 412.76 766.18 417.38 ;
     RECT  780.86 414.86 910.66 417.38 ;
     RECT  921.02 415.28 964.42 417.38 ;
     RECT  1391.9 414.86 1421.38 417.38 ;
     RECT  1433.66 414.02 1444.9 417.38 ;
     RECT  1456.7 414.86 1483.3 417.38 ;
     RECT  1366.94 224.8 1367.14 417.5 ;
     RECT  1511.9 417.38 1512.1 417.5 ;
     RECT  1576.7 397.64 1576.9 417.5 ;
     RECT  1365.98 417.5 1367.14 417.7 ;
     RECT  1576.22 417.5 1576.9 417.7 ;
     RECT  1391.9 417.38 1483.3 417.8 ;
     RECT  1509.98 417.5 1512.1 417.8 ;
     RECT  592.7 415.945 595.78 418.22 ;
     RECT  609.5 415.7 612.58 418.22 ;
     RECT  983.9 416.96 984.58 418.22 ;
     RECT  1528.22 416.54 1559.14 418.22 ;
     RECT  645.98 417.38 766.18 418.64 ;
     RECT  780.86 417.38 967.78 418.64 ;
     RECT  1525.34 418.22 1559.62 418.64 ;
     RECT  460.7 413.6 554.5 419.06 ;
     RECT  566.78 415.945 578.5 419.06 ;
     RECT  592.7 418.22 612.58 419.06 ;
     RECT  622.94 417.8 623.14 419.06 ;
     RECT  645.98 418.64 768.1 419.9 ;
     RECT  780.86 418.64 969.22 419.9 ;
     RECT  645.98 419.9 969.22 420.74 ;
     RECT  981.5 418.22 984.58 420.74 ;
     RECT  1391.9 417.8 1512.1 421.16 ;
     RECT  235.58 416.96 421.06 421.58 ;
     RECT  1386.14 421.16 1512.1 421.58 ;
     RECT  1005.02 415.945 1005.22 422.15 ;
     RECT  1005.02 422.15 1011.52 423.68 ;
     RECT  1386.14 421.58 1512.58 423.68 ;
     RECT  1524.86 418.64 1559.62 423.68 ;
     RECT  1386.14 423.68 1559.62 424.3 ;
     RECT  1386.14 424.3 1558.18 425.56 ;
     RECT  -70 388.4 218.5 427.35 ;
     RECT  229.34 421.58 421.06 427.35 ;
     RECT  437.18 408.56 449.38 427.35 ;
     RECT  459.74 419.06 578.5 427.35 ;
     RECT  592.7 419.06 623.14 427.35 ;
     RECT  645.98 420.74 984.58 427.35 ;
     RECT  994.94 415.945 995.14 427.35 ;
     RECT  1005.02 423.68 1012.42 427.35 ;
     RECT  1331.235 215.315 1336.765 432.08 ;
     RECT  1304.06 432.5 1304.26 432.92 ;
     RECT  1319.42 432.08 1319.62 432.92 ;
     RECT  1331.235 432.08 1340.74 432.92 ;
     RECT  1353.5 432.08 1353.7 432.92 ;
     RECT  1365.98 417.7 1366.18 432.92 ;
     RECT  1295.42 432.92 1304.26 433.34 ;
     RECT  1317.98 432.92 1319.62 433.34 ;
     RECT  1329.5 432.92 1340.74 433.34 ;
     RECT  1351.1 432.92 1366.18 433.34 ;
     RECT  1386.62 425.56 1558.18 435.86 ;
     RECT  1295.42 433.34 1366.18 436.28 ;
     RECT  1381.82 435.86 1558.18 436.28 ;
     RECT  1576.22 417.7 1576.42 436.28 ;
     RECT  1287.26 436.28 1371.46 436.7 ;
     RECT  1284.38 436.7 1371.46 437.54 ;
     RECT  1381.82 436.28 1576.42 437.54 ;
     RECT  -70 427.35 1012.42 439.1 ;
     RECT  1284.38 437.54 1576.42 440.48 ;
     RECT  1281.98 440.48 1576.42 445.94 ;
     RECT  1588.185 381 1870 445.94 ;
     RECT  1260.86 440.48 1261.06 446.78 ;
     RECT  1260.86 446.78 1269.22 447.62 ;
     RECT  1281.98 445.94 1870 447.62 ;
     RECT  -70 439.1 1013.86 451 ;
     RECT  1260.86 447.62 1870 451 ;
     RECT  1260.86 451 1800 451.4 ;
     RECT  1254.62 451.4 1800 455.6 ;
     RECT  0 451 1013.86 469 ;
     RECT  1250.78 455.6 1800 469 ;
     RECT  1250.78 469 1870 474.7 ;
     RECT  1250.78 474.7 1576.42 484.58 ;
     RECT  1588.185 474.7 1870 484.58 ;
     RECT  1250.78 484.58 1870 497.38 ;
     RECT  1251.26 497.38 1870 503.68 ;
     RECT  1251.26 503.68 1576.42 512.08 ;
     RECT  1162.46 507.26 1162.66 518.6 ;
     RECT  1127.235 215.315 1132.765 519.02 ;
     RECT  1155.26 518.6 1162.66 519.02 ;
     RECT  1173.02 518.6 1173.7 519.02 ;
     RECT  1151.9 519.02 1173.7 519.44 ;
     RECT  1195.235 223.96 1200.765 519.44 ;
     RECT  1127.235 519.02 1137.22 519.86 ;
     RECT  1151.9 519.44 1200.765 519.86 ;
     RECT  -70 469 1013.86 520.7 ;
     RECT  1253.18 512.08 1576.42 524.06 ;
     RECT  -70 520.7 1015.3 524.48 ;
     RECT  1127.235 519.86 1200.765 526.58 ;
     RECT  -70 524.48 1018.18 527 ;
     RECT  1253.18 524.06 1577.86 527.2 ;
     RECT  -70 527 1020.58 527.42 ;
     RECT  -70 527.42 1023.94 528.26 ;
     RECT  1253.18 527.2 1576.42 531.2 ;
     RECT  1111.1 531.2 1111.3 531.62 ;
     RECT  1122.62 526.58 1200.765 531.62 ;
     RECT  1111.1 531.62 1200.765 532.88 ;
     RECT  -70 528.26 1030.18 533.08 ;
     RECT  1102.46 532.88 1200.765 534.14 ;
     RECT  1225.82 180 1226.02 534.14 ;
     RECT  1218.14 534.14 1226.02 534.56 ;
     RECT  1102.46 534.14 1202.5 538.76 ;
     RECT  1251.74 531.2 1576.42 538.96 ;
     RECT  -70 533.08 1026.34 539 ;
     RECT  1588.185 503.68 1870 539 ;
     RECT  1095.74 538.76 1202.5 539.38 ;
     RECT  0 539 1026.34 541.9 ;
     RECT  1095.74 539.38 1202.02 543.38 ;
     RECT  0 541.9 1024.9 546.13 ;
     RECT  1036.7 545.9 1053.22 546.32 ;
     RECT  1036.7 546.32 1056.1 548.84 ;
     RECT  1067.42 547.16 1067.62 548.84 ;
     RECT  1036.7 548.84 1071.94 549.26 ;
     RECT  1081.82 546.32 1082.02 549.26 ;
     RECT  1238.3 542.12 1238.5 549.26 ;
     RECT  1255.58 538.96 1576.42 549.26 ;
     RECT  1588.185 539 1800 549.26 ;
     RECT  1036.7 549.26 1082.02 549.68 ;
     RECT  1035.26 549.68 1082.02 550.1 ;
     RECT  1035.26 550.1 1082.5 550.94 ;
     RECT  1093.34 543.38 1202.02 550.94 ;
     RECT  0 546.13 579.94 551.98 ;
     RECT  1237.34 549.26 1238.5 553.04 ;
     RECT  235.58 551.98 579.94 553.24 ;
     RECT  1035.26 550.94 1202.02 553.24 ;
     RECT  1212.86 534.56 1226.02 553.46 ;
     RECT  1237.34 553.04 1245.7 553.46 ;
     RECT  0 551.98 223.78 553.66 ;
     RECT  235.58 553.24 504.58 553.66 ;
     RECT  589.82 546.13 1024.9 553.66 ;
     RECT  847.58 553.66 1024.9 553.88 ;
     RECT  1035.26 553.24 1201.54 553.88 ;
     RECT  1212.86 553.46 1245.7 554.3 ;
     RECT  235.58 553.66 489.22 554.5 ;
     RECT  235.58 554.5 243.94 554.92 ;
     RECT  253.82 554.5 325.06 554.92 ;
     RECT  515.235 553.24 579.94 554.92 ;
     RECT  241.82 554.92 243.94 555.34 ;
     RECT  337.34 554.5 410.5 555.76 ;
     RECT  253.82 554.92 293.38 556.18 ;
     RECT  561.5 554.92 579.94 556.4 ;
     RECT  589.82 553.66 837.22 556.4 ;
     RECT  243.74 555.34 243.94 556.6 ;
     RECT  253.82 556.18 259.3 556.6 ;
     RECT  363.74 555.76 410.5 556.6 ;
     RECT  0 553.66 218.98 557 ;
     RECT  1255.58 549.26 1800 557 ;
     RECT  561.5 556.4 837.22 557.02 ;
     RECT  370.46 556.6 410.5 557.44 ;
     RECT  272.06 556.18 293.38 557.86 ;
     RECT  370.46 557.44 409.06 558.28 ;
     RECT  446.3 554.5 489.22 558.28 ;
     RECT  1211.9 554.3 1245.7 558.5 ;
     RECT  1255.58 557 1870 558.5 ;
     RECT  455.42 558.28 489.22 559.54 ;
     RECT  456.38 559.54 489.22 560.38 ;
     RECT  303.74 554.92 325.06 560.8 ;
     RECT  293.18 557.86 293.38 561.22 ;
     RECT  370.46 558.28 387.94 561.22 ;
     RECT  1211.9 558.5 1870 561.22 ;
     RECT  337.34 555.76 347.62 562.48 ;
     RECT  378.62 561.22 387.94 563.32 ;
     RECT  515.235 554.92 549.7 563.32 ;
     RECT  303.74 560.8 321.7 563.74 ;
     RECT  847.58 553.88 1201.54 564.38 ;
     RECT  1211.9 561.22 1256.74 564.38 ;
     RECT  404.06 558.28 409.06 564.58 ;
     RECT  421.82 554.5 433.06 565 ;
     RECT  404.06 564.58 408.1 565.84 ;
     RECT  456.38 560.38 481.54 566.68 ;
     RECT  561.5 557.02 561.7 567.1 ;
     RECT  303.74 563.74 318.82 568.36 ;
     RECT  378.62 563.32 386.02 568.78 ;
     RECT  572.06 557.02 837.22 569 ;
     RECT  847.58 564.38 1256.74 569 ;
     RECT  -70 557 218.98 573.82 ;
     RECT  255.26 556.6 259.3 574.24 ;
     RECT  421.82 565 428.26 577.18 ;
     RECT  572.06 569 1256.74 578.02 ;
     RECT  500.54 553.66 504.58 578.86 ;
     RECT  583.235 578.02 1256.74 580.34 ;
     RECT  1266.62 561.22 1870 580.34 ;
     RECT  583.235 580.34 1870 584.32 ;
     RECT  311.235 568.36 318.82 588.94 ;
     RECT  748.22 584.32 1870 595.04 ;
     RECT  583.235 584.32 732.1 599.24 ;
     RECT  741.98 595.04 1870 599.24 ;
     RECT  583.235 599.24 1870 599.44 ;
     RECT  428.06 577.18 428.26 600.08 ;
     RECT  379.235 568.78 386.02 601.54 ;
     RECT  456.38 566.68 456.58 602.38 ;
     RECT  583.235 599.44 837.7 602.8 ;
     RECT  583.235 602.8 835.3 603.22 ;
     RECT  583.235 603.22 831.94 604.06 ;
     RECT  583.235 604.06 629.86 604.9 ;
     RECT  583.235 604.9 629.38 606.58 ;
     RECT  272.06 557.86 279.94 608.26 ;
     RECT  583.235 606.58 628.42 608.26 ;
     RECT  404.06 565.84 404.26 609.1 ;
     RECT  473.18 566.68 481.54 609.1 ;
     RECT  850.46 599.44 1870 609.32 ;
     RECT  426.62 600.08 428.26 609.52 ;
     RECT  600.86 608.26 628.42 610.78 ;
     RECT  549.5 563.32 549.7 612.88 ;
     RECT  640.7 604.06 831.94 614.78 ;
     RECT  338.78 562.48 347.62 614.98 ;
     RECT  255.26 574.24 255.46 615.82 ;
     RECT  279.74 608.26 279.94 616.66 ;
     RECT  504.38 578.86 504.58 617.5 ;
     RECT  639.26 614.78 831.94 617.5 ;
     RECT  648.86 617.5 831.94 617.72 ;
     RECT  845.18 609.32 1870 617.72 ;
     RECT  515.235 563.32 527.14 618.56 ;
     RECT  648.86 617.72 1870 619.18 ;
     RECT  338.78 614.98 338.98 619.6 ;
     RECT  572.06 578.02 572.26 621.5 ;
     RECT  648.86 619.18 893.38 621.7 ;
     RECT  649.82 621.7 893.38 622.12 ;
     RECT  654.14 622.12 893.38 622.96 ;
     RECT  508.7 618.56 527.14 623.8 ;
     RECT  555.74 623.18 555.94 624.02 ;
     RECT  311.235 588.94 316.765 624.86 ;
     RECT  379.235 601.54 384.765 625.28 ;
     RECT  237.02 618.98 237.22 625.7 ;
     RECT  655.1 622.96 893.38 626.32 ;
     RECT  481.34 609.1 481.54 626.96 ;
     RECT  -70 573.82 211.815 627 ;
     RECT  903.74 619.18 1870 627 ;
     RECT  481.34 626.96 482.5 627.16 ;
     RECT  600.86 610.78 623.14 627.8 ;
     RECT  415.1 628.64 415.3 629.06 ;
     RECT  406.94 629.06 415.3 630.32 ;
     RECT  426.62 609.52 427.78 630.32 ;
     RECT  311.235 624.86 322.66 630.74 ;
     RECT  571.58 621.5 572.26 631.36 ;
     RECT  309.02 630.74 322.66 631.58 ;
     RECT  600.86 627.8 625.54 631.78 ;
     RECT  839.42 626.32 893.38 631.78 ;
     RECT  237.02 625.7 242.02 633.26 ;
     RECT  279.26 632.84 279.46 633.68 ;
     RECT  237.02 633.26 242.98 634.1 ;
     RECT  583.235 608.26 588.765 634.94 ;
     RECT  399.74 630.32 427.78 635.36 ;
     RECT  655.1 626.32 829.54 636.2 ;
     RECT  839.42 631.78 873.22 636.2 ;
     RECT  544.22 635.78 544.42 636.62 ;
     RECT  508.7 623.8 520.765 637.04 ;
     RECT  655.1 636.2 873.22 637.04 ;
     RECT  903.74 627 1800 637.24 ;
     RECT  370.46 625.28 384.765 637.46 ;
     RECT  399.74 635.36 432.58 637.46 ;
     RECT  583.235 634.94 590.02 637.88 ;
     RECT  600.86 631.78 602.02 637.88 ;
     RECT  651.74 637.04 873.22 637.88 ;
     RECT  302.78 631.58 322.66 638.72 ;
     RECT  887.42 631.78 893.38 638.72 ;
     RECT  903.74 637.24 960.58 638.72 ;
     RECT  302.78 638.72 325.06 639.14 ;
     RECT  370.46 637.46 432.58 640.7 ;
     RECT  466.94 639.56 467.14 640.82 ;
     RECT  482.3 627.16 482.5 640.82 ;
     RECT  571.58 631.36 571.78 641.24 ;
     RECT  583.235 637.88 602.02 641.24 ;
     RECT  466.94 640.82 482.5 641.66 ;
     RECT  445.82 629.48 446.02 642.5 ;
     RECT  614.78 631.78 625.54 643.34 ;
     RECT  0 627 211.815 645 ;
     RECT  970.46 637.24 1800 645 ;
     RECT  649.82 637.88 873.22 645.02 ;
     RECT  300.38 639.14 325.06 645.44 ;
     RECT  343.1 632.42 343.3 645.86 ;
     RECT  355.58 632 355.78 645.86 ;
     RECT  648.38 645.02 877.54 645.86 ;
     RECT  887.42 638.72 960.58 645.86 ;
     RECT  279.26 633.68 281.38 646.7 ;
     RECT  297.02 645.44 325.06 646.7 ;
     RECT  445.82 642.5 455.14 646.7 ;
     RECT  465.98 641.66 482.5 646.7 ;
     RECT  237.02 634.1 243.46 647.12 ;
     RECT  224.06 634.52 224.26 647.54 ;
     RECT  235.1 647.12 243.46 647.54 ;
     RECT  279.26 646.7 325.06 648.38 ;
     RECT  648.38 645.86 960.58 648.38 ;
     RECT  970.46 645 1870 648.38 ;
     RECT  571.58 641.24 602.02 648.8 ;
     RECT  555.74 624.02 556.9 650.9 ;
     RECT  648.38 648.38 1870 652.16 ;
     RECT  370.46 640.7 433.54 652.58 ;
     RECT  343.1 645.86 355.78 653 ;
     RECT  367.1 652.58 433.54 653 ;
     RECT  640.7 652.16 1870 653.2 ;
     RECT  343.1 653 433.54 653.84 ;
     RECT  501.02 637.04 520.765 655.1 ;
     RECT  555.74 650.9 560.74 655.52 ;
     RECT  614.78 643.34 628.42 655.52 ;
     RECT  542.3 636.62 545.38 656.36 ;
     RECT  224.06 647.54 243.46 656.78 ;
     RECT  614.78 655.52 629.86 656.78 ;
     RECT  445.82 646.7 482.5 657.2 ;
     RECT  495.26 655.1 520.765 657.2 ;
     RECT  555.74 655.52 561.7 658.04 ;
     RECT  571.58 648.8 603.46 658.04 ;
     RECT  336.38 653.84 433.54 658.46 ;
     RECT  445.82 657.2 520.765 658.46 ;
     RECT  336.38 658.46 520.765 660.56 ;
     RECT  535.1 656.36 545.38 660.56 ;
     RECT  224.06 656.78 243.94 663.08 ;
     RECT  648.38 653.2 1870 663.28 ;
     RECT  336.38 660.56 545.38 663.5 ;
     RECT  555.74 658.04 603.46 663.5 ;
     RECT  614.78 656.78 630.34 663.92 ;
     RECT  648.38 663.28 1053.7 665.6 ;
     RECT  272.54 648.38 325.06 666.02 ;
     RECT  1063.58 663.28 1870 667.48 ;
     RECT  647.42 665.6 1053.7 667.7 ;
     RECT  646.94 667.7 1053.7 668.12 ;
     RECT  614.78 663.92 636.58 668.96 ;
     RECT  646.46 668.12 1053.7 668.96 ;
     RECT  614.78 668.96 1053.7 669.8 ;
     RECT  1318.94 667.48 1870 672.52 ;
     RECT  336.38 663.5 603.46 672.74 ;
     RECT  613.34 669.8 1053.7 672.74 ;
     RECT  336.38 672.74 1053.7 674 ;
     RECT  1063.58 667.48 1305.7 674 ;
     RECT  224.06 663.08 248.26 675.68 ;
     RECT  224.06 675.68 257.86 676.1 ;
     RECT  271.58 666.02 325.06 676.1 ;
     RECT  336.38 674 1305.7 682.82 ;
     RECT  1319.9 672.52 1870 682.82 ;
     RECT  224.06 676.1 325.06 684.92 ;
     RECT  336.38 682.82 1870 684.92 ;
     RECT  224.06 684.92 1870 690.16 ;
     RECT  -70 645 211.815 698.36 ;
     RECT  224.06 690.16 627.46 698.36 ;
     RECT  -70 698.36 627.46 702.98 ;
     RECT  639.74 690.16 1870 705.28 ;
     RECT  -70 702.98 628.42 709.25 ;
     RECT  639.74 705.28 1310.02 709.25 ;
     RECT  -70 709.25 1310.02 715 ;
     RECT  1323.26 705.28 1870 715 ;
     RECT  0 715 1310.02 716 ;
     RECT  1323.26 715 1800 716 ;
     RECT  0 716 1800 733 ;
     RECT  -70 733 1870 735.1 ;
     RECT  -70 735.1 1578.34 743.08 ;
     RECT  -70 743.08 1472.26 745.6 ;
     RECT  1486.46 743.08 1578.34 746.02 ;
     RECT  1497.98 746.02 1578.34 746.86 ;
     RECT  -70 745.6 1470.82 750.64 ;
     RECT  1498.46 746.86 1561.06 750.64 ;
     RECT  1524.38 750.64 1546.66 751.06 ;
     RECT  1560.86 750.64 1561.06 751.06 ;
     RECT  1498.46 750.64 1514.02 753.58 ;
     RECT  1529.66 751.06 1546.66 753.58 ;
     RECT  1498.46 753.58 1511.14 754 ;
     RECT  1530.14 753.58 1546.66 754 ;
     RECT  1499.9 754 1511.14 754.84 ;
     RECT  1530.62 754 1546.66 754.84 ;
     RECT  1501.34 754.84 1511.14 756.52 ;
     RECT  1501.34 756.52 1504.9 757.36 ;
     RECT  -70 750.64 1466.98 770.38 ;
     RECT  1486.46 746.02 1486.66 775.42 ;
     RECT  1501.34 757.36 1504.42 781.1 ;
     RECT  -70 770.38 1457.38 787.6 ;
     RECT  1497.02 781.1 1504.42 788.44 ;
     RECT  1468.7 775.22 1468.9 802.3 ;
     RECT  -70 787.6 1454.5 803 ;
     RECT  1588.185 735.1 1870 803 ;
     RECT  1558.46 802.52 1558.66 807.98 ;
     RECT  1574.3 746.86 1578.34 807.98 ;
     RECT  0 803 1454.5 821 ;
     RECT  1588.185 803 1800 821 ;
     RECT  1558.46 807.98 1578.34 821.62 ;
     RECT  -70 821 1454.5 828.03 ;
     RECT  -70 828.03 217.64 830.63 ;
     RECT  655.1 828.03 1454.5 832.76 ;
     RECT  -70 830.63 215.04 833.23 ;
     RECT  334.46 828.03 334.66 833.8 ;
     RECT  655.1 832.76 1455.94 834.44 ;
     RECT  1558.46 821.62 1576.9 837.8 ;
     RECT  593.66 828.03 593.86 839.015 ;
     RECT  583.235 839.015 593.86 840.74 ;
     RECT  553.82 841.16 554.02 842 ;
     RECT  583.235 840.74 594.82 842 ;
     RECT  640.22 828.03 640.42 842 ;
     RECT  655.1 834.44 1463.62 842 ;
     RECT  546.62 842 554.02 847.88 ;
     RECT  515.235 828.03 520.765 848.3 ;
     RECT  623.42 849.56 623.62 849.98 ;
     RECT  640.22 842 1463.62 849.98 ;
     RECT  565.82 839.9 566.02 851.24 ;
     RECT  501.02 853.76 501.22 854.6 ;
     RECT  481.82 852.08 482.02 855.86 ;
     RECT  277.82 855.86 278.02 856.28 ;
     RECT  277.82 856.28 280.9 856.7 ;
     RECT  240.86 828.03 242.98 857.54 ;
     RECT  583.235 842 597.22 857.96 ;
     RECT  611.42 849.14 611.62 857.96 ;
     RECT  501.02 854.6 503.62 858.38 ;
     RECT  515.235 848.3 522.82 858.38 ;
     RECT  277.82 856.7 281.86 859.64 ;
     RECT  276.38 859.64 281.86 860.06 ;
     RECT  438.62 859.22 438.82 860.9 ;
     RECT  501.02 858.38 522.82 862.16 ;
     RECT  537.02 847.88 554.02 862.16 ;
     RECT  477.02 855.86 482.02 862.58 ;
     RECT  263.42 863 263.62 863.84 ;
     RECT  276.38 860.06 282.82 863.84 ;
     RECT  295.1 863 295.3 863.84 ;
     RECT  1558.46 837.8 1578.34 864.04 ;
     RECT  472.22 862.58 482.02 864.68 ;
     RECT  263.42 863.84 295.3 866.98 ;
     RECT  565.82 851.24 570.82 867.2 ;
     RECT  583.235 857.96 611.62 867.2 ;
     RECT  269.18 866.98 295.3 867.4 ;
     RECT  269.18 867.4 283.78 868.24 ;
     RECT  501.02 862.16 554.02 868.46 ;
     RECT  235.58 857.54 242.98 869.72 ;
     RECT  269.18 868.24 279.94 870.34 ;
     RECT  235.58 869.72 244.9 870.98 ;
     RECT  472.22 864.68 484.42 870.98 ;
     RECT  565.82 867.2 611.62 870.98 ;
     RECT  623.42 849.98 1463.62 870.98 ;
     RECT  294.62 867.4 295.3 871.6 ;
     RECT  498.62 868.46 554.02 871.82 ;
     RECT  269.18 870.34 278.02 872.02 ;
     RECT  277.82 872.02 278.02 872.86 ;
     RECT  296.54 872.24 296.74 872.86 ;
     RECT  311.235 828.03 316.765 873.325 ;
     RECT  465.02 870.98 484.42 873.5 ;
     RECT  496.22 871.82 554.02 873.5 ;
     RECT  465.02 873.5 554.02 874.76 ;
     RECT  565.82 870.98 1463.62 874.76 ;
     RECT  -70 833.23 211.815 875.6 ;
     RECT  438.62 860.9 446.02 875.6 ;
     RECT  438.62 875.6 450.82 876.02 ;
     RECT  465.02 874.76 1463.62 876.02 ;
     RECT  379.235 839.015 384.765 877.105 ;
     RECT  438.62 876.02 1463.62 878.96 ;
     RECT  438.62 878.96 1464.58 880.88 ;
     RECT  441.02 880.88 1464.58 881.3 ;
     RECT  443.42 881.3 1464.58 882.14 ;
     RECT  445.82 882.14 1464.58 882.98 ;
     RECT  510.62 882.98 1464.58 883.4 ;
     RECT  769.82 883.4 1464.58 883.58 ;
     RECT  510.62 883.4 755.62 883.82 ;
     RECT  445.82 882.98 498.82 884.24 ;
     RECT  445.82 884.24 496.42 884.66 ;
     RECT  445.82 884.66 491.62 885.5 ;
     RECT  510.62 883.82 570.82 887.18 ;
     RECT  587.42 883.82 755.62 887.6 ;
     RECT  769.82 883.58 1467.46 889.04 ;
     RECT  1535.235 754.84 1546.66 889.04 ;
     RECT  769.82 889.04 1467.94 889.88 ;
     RECT  727.1 887.6 755.62 890.12 ;
     RECT  -70 875.6 216.1 891 ;
     RECT  1588.185 821 1870 891 ;
     RECT  510.62 887.18 566.02 891.38 ;
     RECT  1497.02 788.44 1497.22 892.7 ;
     RECT  1496.54 892.7 1497.22 892.9 ;
     RECT  769.82 889.88 1468.9 893.44 ;
     RECT  610.94 887.6 668.74 894.32 ;
     RECT  727.1 890.12 753.22 897.68 ;
     RECT  769.82 893.44 1467.94 901.42 ;
     RECT  612.38 894.32 668.74 903.78 ;
     RECT  678.62 887.6 715.78 903.78 ;
     RECT  727.1 897.68 746.02 903.78 ;
     RECT  769.82 901.42 1467.46 903.78 ;
     RECT  587.42 887.6 594.34 904.62 ;
     RECT  612.38 903.78 746.02 904.62 ;
     RECT  765.5 903.78 1467.46 905.04 ;
     RECT  587.42 904.62 746.02 906.72 ;
     RECT  370.94 907.14 371.14 907.56 ;
     RECT  445.82 885.5 484.42 907.56 ;
     RECT  510.62 891.38 540.58 907.56 ;
     RECT  350.3 907.56 350.5 907.98 ;
     RECT  370.94 907.56 377.86 907.98 ;
     RECT  441.02 907.56 484.42 907.98 ;
     RECT  503.9 907.56 540.58 907.98 ;
     RECT  551.42 891.38 566.02 907.98 ;
     RECT  579.74 906.72 746.02 907.98 ;
     RECT  756.38 905.04 1467.46 907.98 ;
     RECT  414.14 907.56 414.34 908.4 ;
     RECT  430.46 906.3 430.66 908.4 ;
     RECT  441.02 907.98 1467.46 908.4 ;
     RECT  394.94 908.4 395.14 908.82 ;
     RECT  408.38 908.4 414.34 908.82 ;
     RECT  0 891 216.1 909 ;
     RECT  1588.185 891 1800 909 ;
     RECT  349.82 907.98 350.5 909.24 ;
     RECT  360.86 907.98 379.78 909.24 ;
     RECT  394.94 908.82 414.34 910.5 ;
     RECT  394.46 910.5 414.34 910.92 ;
     RECT  424.22 908.4 1467.46 910.92 ;
     RECT  349.82 909.24 379.78 911.34 ;
     RECT  394.46 910.92 1467.46 911.72 ;
     RECT  394.46 911.72 1472.74 912.56 ;
     RECT  349.82 911.34 384.1 912.6 ;
     RECT  394.46 912.56 1473.22 912.6 ;
     RECT  349.82 912.6 1473.22 914.66 ;
     RECT  349.82 914.66 1481.38 915.12 ;
     RECT  349.34 915.12 1481.38 915.54 ;
     RECT  345.5 915.54 1481.38 915.92 ;
     RECT  334.46 915.12 335.14 915.96 ;
     RECT  333.98 915.96 335.14 916.38 ;
     RECT  345.5 915.92 1482.34 916.38 ;
     RECT  333.98 916.38 1482.34 918.9 ;
     RECT  333.02 918.9 1482.34 919.32 ;
     RECT  329.66 919.32 1482.34 920.12 ;
     RECT  1496.54 892.9 1496.74 920.12 ;
     RECT  329.66 920.12 1496.74 920.54 ;
     RECT  319.1 918.9 319.3 923.1 ;
     RECT  315.26 923.1 319.3 923.94 ;
     RECT  329.66 920.54 1504.9 923.94 ;
     RECT  1565.66 864.04 1578.34 925.58 ;
     RECT  1588.185 909 1870 925.58 ;
     RECT  311.42 923.94 1504.9 926.84 ;
     RECT  1565.66 925.58 1870 928.94 ;
     RECT  1558.46 928.94 1870 929.14 ;
     RECT  311.42 926.84 1511.14 930.44 ;
     RECT  312.38 930.44 1511.14 942.8 ;
     RECT  312.38 942.8 1511.62 942.84 ;
     RECT  235.58 870.98 245.38 944.06 ;
     RECT  306.14 942.84 1511.62 945.78 ;
     RECT  302.3 945.78 1511.62 951.62 ;
     RECT  302.3 951.62 1512.1 952.92 ;
     RECT  298.94 952.92 1512.1 956.28 ;
     RECT  291.74 956.28 1512.1 962.12 ;
     RECT  1529.66 889.04 1546.66 964.84 ;
     RECT  277.34 964.26 277.54 965.1 ;
     RECT  291.74 962.12 1515.94 965.1 ;
     RECT  277.34 965.1 1515.94 968.46 ;
     RECT  271.58 968.46 1515.94 969.68 ;
     RECT  271.58 969.68 1519.78 971.4 ;
     RECT  1535.235 964.84 1546.66 972.2 ;
     RECT  1558.46 929.14 1558.66 972.2 ;
     RECT  1535.235 972.2 1558.66 972.4 ;
     RECT  262.94 971.4 1519.78 974.5 ;
     RECT  262.94 974.5 1519.3 974.96 ;
     RECT  -70 909 216.1 979 ;
     RECT  1574.3 929.14 1870 979 ;
     RECT  1574.3 979 1800 979.34 ;
     RECT  264.86 974.96 1519.3 980.8 ;
     RECT  264.86 980.8 1517.38 986.94 ;
     RECT  262.94 986.94 1517.38 988.36 ;
     RECT  1494.14 988.36 1517.38 989.2 ;
     RECT  262.94 988.36 1484.26 990.3 ;
     RECT  1494.14 989.2 1514.5 992.14 ;
     RECT  233.66 944.06 245.38 994.5 ;
     RECT  260.06 990.3 1484.26 994.5 ;
     RECT  1496.54 992.14 1514.5 994.66 ;
     RECT  233.66 994.5 1484.26 995.08 ;
     RECT  1496.54 994.66 1508.74 995.92 ;
     RECT  1496.54 995.92 1505.86 996.34 ;
     RECT  0 979 216.1 997 ;
     RECT  1572.86 979.34 1800 997 ;
     RECT  233.66 995.08 1483.3 1003.48 ;
     RECT  1315.58 1003.48 1483.3 1009.16 ;
     RECT  1315.58 1009.16 1486.66 1010.84 ;
     RECT  1496.54 996.34 1496.74 1010.84 ;
     RECT  233.66 1003.48 1305.7 1011.04 ;
     RECT  1292.06 1011.04 1305.7 1015.04 ;
     RECT  1315.58 1010.84 1497.22 1015.04 ;
     RECT  1292.06 1015.04 1497.22 1015.24 ;
     RECT  1303.1 1015.24 1497.22 1027.42 ;
     RECT  1535.235 972.4 1551.94 1029.52 ;
     RECT  233.66 1011.04 1282.18 1030.36 ;
     RECT  233.66 1030.36 1280.26 1037.12 ;
     RECT  1303.1 1027.42 1373.38 1037.3 ;
     RECT  1383.74 1027.42 1497.22 1037.3 ;
     RECT  888.38 1037.12 1280.26 1041.5 ;
     RECT  1292.06 1015.24 1292.26 1041.5 ;
     RECT  1303.1 1037.3 1497.22 1044.22 ;
     RECT  1303.1 1044.22 1307.14 1044.64 ;
     RECT  1320.38 1044.22 1497.22 1045.28 ;
     RECT  1320.38 1045.28 1498.18 1045.48 ;
     RECT  233.66 1037.12 878.02 1046.78 ;
     RECT  233.66 1046.78 865.54 1047.2 ;
     RECT  1322.3 1045.48 1497.7 1048.84 ;
     RECT  233.66 1047.2 863.14 1049.72 ;
     RECT  888.38 1041.5 1292.26 1050.1 ;
     RECT  1322.3 1048.84 1492.42 1051.78 ;
     RECT  1322.3 1051.78 1489.06 1052.62 ;
     RECT  1322.3 1052.62 1478.02 1053.46 ;
     RECT  1065.5 1050.1 1292.26 1054.94 ;
     RECT  1488.38 1052.62 1489.06 1055.56 ;
     RECT  1322.3 1053.46 1352.74 1056.4 ;
     RECT  1488.38 1055.56 1488.58 1056.4 ;
     RECT  1535.235 1029.52 1551.46 1058.3 ;
     RECT  233.66 1049.72 862.18 1059.38 ;
     RECT  847.1 1059.38 862.18 1060.52 ;
     RECT  847.1 1060.52 861.7 1061.06 ;
     RECT  233.66 1059.38 833.86 1061.9 ;
     RECT  233.66 1061.9 830.02 1062.74 ;
     RECT  233.66 1062.74 829.06 1063.16 ;
     RECT  850.94 1061.06 861.7 1063.58 ;
     RECT  888.38 1050.1 1055.14 1063.76 ;
     RECT  1065.5 1054.94 1295.14 1063.76 ;
     RECT  1323.74 1056.4 1352.74 1063.76 ;
     RECT  1364.54 1053.46 1478.02 1063.76 ;
     RECT  1572.86 997 1870 1065.44 ;
     RECT  -70 997 216.1 1067 ;
     RECT  1565.66 1065.44 1870 1067 ;
     RECT  1491.74 1066.7 1491.94 1067.12 ;
     RECT  1491.74 1067.12 1499.14 1067.54 ;
     RECT  1323.74 1063.76 1478.02 1068.8 ;
     RECT  1491.74 1067.54 1507.78 1068.8 ;
     RECT  1323.74 1068.8 1507.78 1071.74 ;
     RECT  233.66 1063.16 820.9 1074.3 ;
     RECT  1306.94 1044.64 1307.14 1074.68 ;
     RECT  1323.74 1071.74 1512.1 1074.68 ;
     RECT  1306.94 1074.68 1512.1 1075.94 ;
     RECT  888.38 1063.76 1295.14 1078.46 ;
     RECT  1306.94 1075.94 1520.74 1078.46 ;
     RECT  233.66 1074.3 824.74 1082.7 ;
     RECT  233.66 1082.7 827.14 1083.12 ;
     RECT  850.94 1063.58 858.34 1084.58 ;
     RECT  0 1067 216.1 1085 ;
     RECT  1565.66 1067 1800 1085 ;
     RECT  233.66 1083.12 831.46 1085.22 ;
     RECT  856.22 1084.58 858.34 1087.1 ;
     RECT  888.38 1078.46 1520.74 1091.48 ;
     RECT  1534.46 1058.3 1551.46 1091.48 ;
     RECT  233.66 1085.22 831.94 1092.78 ;
     RECT  233.66 1092.78 838.66 1096.76 ;
     RECT  888.38 1091.48 1551.46 1099.66 ;
     RECT  233.66 1096.76 833.38 1111.46 ;
     RECT  233.66 1111.46 832.9 1111.88 ;
     RECT  1551.26 1099.66 1551.46 1115.84 ;
     RECT  888.38 1099.66 1540.765 1116.04 ;
     RECT  1565.66 1085 1870 1116.04 ;
     RECT  -70 1085 216.1 1118.78 ;
     RECT  1535.235 1116.04 1540.765 1119.62 ;
     RECT  1551.26 1115.84 1555.3 1119.62 ;
     RECT  1573.82 1116.04 1870 1119.82 ;
     RECT  233.66 1111.88 831.94 1121.54 ;
     RECT  233.66 1121.54 829.54 1122.38 ;
     RECT  233.66 1122.38 827.14 1127 ;
     RECT  888.38 1116.04 1525.54 1128.44 ;
     RECT  1535.235 1119.62 1555.3 1128.44 ;
     RECT  233.66 1127 824.74 1129.94 ;
     RECT  233.66 1129.94 817.06 1130.36 ;
     RECT  233.66 1130.36 816.58 1130.78 ;
     RECT  233.66 1130.78 571.3 1132.46 ;
     RECT  582.14 1130.78 816.58 1133.72 ;
     RECT  583.1 1133.72 816.58 1134.56 ;
     RECT  553.82 1132.46 571.3 1134.98 ;
     RECT  583.1 1134.56 811.3 1134.98 ;
     RECT  233.66 1132.46 543.46 1135.4 ;
     RECT  583.1 1134.98 583.3 1135.4 ;
     RECT  783.74 1134.98 785.38 1135.4 ;
     RECT  799.1 1134.98 806.5 1135.4 ;
     RECT  785.18 1135.4 785.38 1136.24 ;
     RECT  877.82 1046.78 878.02 1136.42 ;
     RECT  888.38 1128.44 1555.3 1136.42 ;
     RECT  594.14 1134.98 770.5 1136.66 ;
     RECT  556.22 1134.98 564.58 1137.08 ;
     RECT  556.22 1137.08 556.42 1137.5 ;
     RECT  599.9 1136.66 770.5 1137.5 ;
     RECT  599.9 1137.5 766.18 1142.12 ;
     RECT  233.66 1135.4 537.7 1143.38 ;
     RECT  877.82 1136.42 1555.3 1144.6 ;
     RECT  233.66 1143.38 536.26 1149.68 ;
     RECT  561.02 1152.04 561.22 1153.3 ;
     RECT  561.02 1153.3 563.62 1153.72 ;
     RECT  776.06 1153.3 776.26 1153.72 ;
     RECT  806.3 1135.4 806.5 1154.14 ;
     RECT  586.46 1151.62 586.66 1154.98 ;
     RECT  603.26 1142.12 766.18 1154.98 ;
     RECT  -70 1118.78 219.46 1155 ;
     RECT  1588.185 1119.82 1870 1155 ;
     RECT  586.46 1154.98 766.18 1157.08 ;
     RECT  822.62 1154.56 822.82 1157.08 ;
     RECT  833.66 1137.76 833.86 1157.08 ;
     RECT  561.02 1153.72 567.46 1158.76 ;
     RECT  579.26 1157.08 766.18 1160.44 ;
     RECT  776.06 1153.72 780.1 1160.44 ;
     RECT  512.54 1149.68 536.26 1161.12 ;
     RECT  556.22 1158.76 567.46 1161.28 ;
     RECT  822.62 1157.08 833.86 1161.7 ;
     RECT  579.26 1160.44 780.1 1163.8 ;
     RECT  551.42 1161.28 567.46 1164.22 ;
     RECT  551.42 1164.22 568.42 1164.64 ;
     RECT  578.78 1163.8 780.1 1164.64 ;
     RECT  512.06 1161.12 536.26 1167.16 ;
     RECT  512.06 1167.16 538.66 1167.58 ;
     RECT  551.42 1164.64 780.1 1167.58 ;
     RECT  233.66 1149.68 502.18 1169.26 ;
     RECT  512.06 1167.58 780.1 1169.26 ;
     RECT  0 1155 219.46 1173 ;
     RECT  1588.185 1155 1800 1173 ;
     RECT  804.86 1154.14 806.5 1173.46 ;
     RECT  233.66 1169.26 780.1 1173.88 ;
     RECT  233.66 1173.88 786.34 1174.3 ;
     RECT  801.02 1173.46 806.5 1174.3 ;
     RECT  822.62 1161.7 841.54 1174.3 ;
     RECT  877.82 1144.6 1551.46 1175.14 ;
     RECT  233.66 1174.3 808.42 1175.56 ;
     RECT  818.3 1174.3 841.54 1175.56 ;
     RECT  233.66 1175.56 841.54 1176.82 ;
     RECT  1573.82 1119.82 1578.34 1177.16 ;
     RECT  233.66 1176.82 843.94 1178.08 ;
     RECT  856.22 1087.1 856.42 1178.08 ;
     RECT  868.7 1175.14 1551.46 1178.08 ;
     RECT  233.66 1178.08 1551.46 1181.36 ;
     RECT  1573.34 1177.16 1578.34 1184.72 ;
     RECT  1572.86 1184.72 1578.34 1189.76 ;
     RECT  1588.185 1173 1870 1189.76 ;
     RECT  1572.86 1189.76 1870 1190.38 ;
     RECT  233.66 1181.36 1553.38 1192.9 ;
     RECT  -70 1173 219.46 1243 ;
     RECT  1573.34 1190.38 1870 1243 ;
     RECT  233.66 1192.9 1551.46 1249.6 ;
     RECT  233.66 1249.6 1228.42 1260.32 ;
     RECT  233.66 1260.32 1231.78 1260.74 ;
     RECT  1241.66 1249.6 1551.46 1260.74 ;
     RECT  0 1243 219.46 1261 ;
     RECT  1573.34 1243 1800 1261 ;
     RECT  233.66 1260.74 1551.46 1261.36 ;
     RECT  1573.34 1261 1870 1264.52 ;
     RECT  1252.7 1261.36 1551.46 1271.02 ;
     RECT  1252.7 1271.02 1544.26 1272.28 ;
     RECT  1569.5 1264.52 1870 1274.6 ;
     RECT  233.66 1261.36 1241.86 1276.7 ;
     RECT  1256.54 1272.28 1544.26 1279.84 ;
     RECT  1565.66 1274.6 1870 1285.3 ;
     RECT  233.66 1276.7 1244.74 1288.66 ;
     RECT  1259.9 1279.84 1544.26 1291.6 ;
     RECT  233.66 1288.66 1241.38 1293.28 ;
     RECT  1569.5 1285.3 1870 1293.28 ;
     RECT  903.26 1293.28 1241.38 1294.96 ;
     RECT  1573.34 1293.28 1870 1294.96 ;
     RECT  1261.82 1291.6 1544.26 1302.1 ;
     RECT  1265.18 1302.1 1544.26 1305.88 ;
     RECT  233.66 1293.28 888.58 1307.78 ;
     RECT  903.26 1294.96 1236.1 1307.78 ;
     RECT  1265.66 1305.88 1523.14 1308.82 ;
     RECT  1265.66 1308.82 1460.26 1310.08 ;
     RECT  1267.1 1310.08 1454.98 1313.02 ;
     RECT  1267.1 1313.02 1312.42 1313.44 ;
     RECT  1269.98 1313.44 1312.42 1313.86 ;
     RECT  1269.98 1313.86 1275.94 1314.28 ;
     RECT  1286.78 1313.86 1312.42 1314.28 ;
     RECT  1305.02 1314.28 1312.42 1316.38 ;
     RECT  1286.78 1314.28 1289.38 1317.64 ;
     RECT  1309.82 1316.38 1312.42 1318.06 ;
     RECT  1309.82 1318.06 1310.02 1318.9 ;
     RECT  233.66 1307.78 1236.1 1319.32 ;
     RECT  1470.62 1308.82 1523.14 1321 ;
     RECT  1522.94 1321 1523.14 1321.42 ;
     RECT  1471.58 1321 1505.86 1321.84 ;
     RECT  1323.26 1313.02 1454.98 1322.06 ;
     RECT  1471.58 1321.84 1482.34 1322.26 ;
     RECT  1323.26 1322.06 1456.9 1323.94 ;
     RECT  1288.7 1317.64 1289.38 1324.78 ;
     RECT  1323.26 1323.94 1382.98 1324.78 ;
     RECT  1471.58 1322.26 1479.46 1324.78 ;
     RECT  233.66 1319.32 904.9 1324.82 ;
     RECT  1367.9 1324.78 1382.5 1325.2 ;
     RECT  1477.34 1324.78 1479.46 1325.2 ;
     RECT  1496.54 1321.84 1505.86 1325.2 ;
     RECT  1323.26 1324.78 1357.06 1325.62 ;
     RECT  1575.74 1294.96 1870 1325.84 ;
     RECT  1288.7 1324.78 1288.9 1326.46 ;
     RECT  233.66 1324.82 252.1 1327.34 ;
     RECT  1325.18 1325.62 1357.06 1327.72 ;
     RECT  1392.86 1323.94 1451.14 1327.72 ;
     RECT  1434.62 1327.72 1436.74 1328.14 ;
     RECT  1535.235 1305.88 1544.26 1328.36 ;
     RECT  1325.18 1327.72 1346.98 1328.56 ;
     RECT  1368.38 1325.2 1382.5 1328.56 ;
     RECT  1392.86 1327.72 1420.9 1328.56 ;
     RECT  1435.1 1328.14 1436.74 1328.56 ;
     RECT  1326.14 1328.56 1346.98 1328.98 ;
     RECT  1435.58 1328.56 1436.74 1328.98 ;
     RECT  914.78 1319.32 1236.1 1329.62 ;
     RECT  1392.86 1328.56 1419.46 1330.24 ;
     RECT  262.94 1324.82 904.9 1330.88 ;
     RECT  914.78 1329.62 1238.5 1330.88 ;
     RECT  -70 1261 219.46 1331 ;
     RECT  1574.78 1325.84 1870 1331 ;
     RECT  1392.86 1330.24 1414.18 1331.92 ;
     RECT  1436.54 1328.98 1436.74 1331.92 ;
     RECT  262.94 1330.88 1238.5 1331.96 ;
     RECT  1326.14 1328.98 1340.26 1332.34 ;
     RECT  1326.14 1332.34 1336.765 1332.76 ;
     RECT  1370.78 1328.56 1382.02 1332.76 ;
     RECT  1392.86 1331.92 1410.82 1332.76 ;
     RECT  1450.94 1327.72 1451.14 1332.76 ;
     RECT  1392.86 1332.76 1404.765 1333.6 ;
     RECT  1533.5 1328.36 1544.26 1333.6 ;
     RECT  264.38 1331.96 1238.5 1334.48 ;
     RECT  1535.235 1333.6 1544.26 1334.86 ;
     RECT  266.3 1334.48 1238.5 1336.12 ;
     RECT  1574.78 1331 1800 1339.9 ;
     RECT  266.3 1336.12 1237.54 1340.32 ;
     RECT  1574.78 1339.9 1576.9 1340.32 ;
     RECT  266.3 1340.32 1235.62 1342.04 ;
     RECT  289.82 1342.04 1235.62 1342.46 ;
     RECT  266.3 1342.04 278.98 1343.3 ;
     RECT  278.78 1343.3 278.98 1346.66 ;
     RECT  289.82 1342.46 294.34 1346.66 ;
     RECT  289.82 1346.66 290.02 1347.08 ;
     RECT  306.62 1342.46 1235.62 1347.88 ;
     RECT  0 1331 219.46 1349 ;
     RECT  1588.185 1339.9 1800 1349 ;
     RECT  1221.98 1347.88 1235.62 1354.18 ;
     RECT  1574.78 1340.32 1575.94 1354.4 ;
     RECT  1535.235 1334.86 1540.765 1354.82 ;
     RECT  1221.98 1354.18 1232.26 1355.02 ;
     RECT  1222.94 1355.02 1232.26 1355.44 ;
     RECT  1362.62 1355.66 1362.82 1356.08 ;
     RECT  306.62 1347.88 1210.18 1357.58 ;
     RECT  327.26 1357.58 1210.18 1358 ;
     RECT  338.78 1358 1210.18 1358.6 ;
     RECT  266.3 1343.3 266.5 1359.26 ;
     RECT  1526.3 1354.82 1540.765 1360.7 ;
     RECT  1526.3 1360.7 1547.62 1360.9 ;
     RECT  327.26 1358 327.94 1362.62 ;
     RECT  1357.34 1356.08 1362.82 1363 ;
     RECT  1362.62 1363 1362.82 1363.22 ;
     RECT  1222.94 1355.44 1223.14 1363.42 ;
     RECT  338.78 1358.6 1211.14 1364.26 ;
     RECT  338.78 1364.26 1210.18 1364.3 ;
     RECT  327.26 1362.62 327.46 1364.72 ;
     RECT  306.62 1357.58 314.98 1367.66 ;
     RECT  339.26 1364.3 1210.18 1368.04 ;
     RECT  314.78 1367.66 314.98 1369.34 ;
     RECT  339.26 1368.04 1067.14 1370.56 ;
     RECT  1077.02 1368.04 1210.18 1371.4 ;
     RECT  1535.235 1360.9 1547.62 1378.76 ;
     RECT  1574.78 1354.4 1576.9 1378.76 ;
     RECT  1077.5 1371.4 1210.18 1378.96 ;
     RECT  1535.235 1378.76 1548.1 1378.96 ;
     RECT  339.26 1370.56 1051.3 1380.26 ;
     RECT  1077.5 1378.96 1144.9 1381.48 ;
     RECT  341.66 1380.26 1051.3 1382.12 ;
     RECT  1062.14 1370.56 1062.34 1382.12 ;
     RECT  341.66 1382.12 1062.34 1384.46 ;
     RECT  1159.1 1378.96 1210.18 1385.26 ;
     RECT  1164.86 1385.26 1210.18 1385.68 ;
     RECT  1569.5 1378.76 1576.9 1385.68 ;
     RECT  346.94 1384.46 1062.34 1385.76 ;
     RECT  1399.235 1333.6 1404.765 1386.32 ;
     RECT  492.86 1385.76 1062.34 1388.42 ;
     RECT  1077.5 1381.48 1140.1 1390.1 ;
     RECT  346.94 1385.76 482.5 1390.76 ;
     RECT  346.94 1390.76 477.22 1391.6 ;
     RECT  1074.14 1390.1 1140.1 1391.98 ;
     RECT  492.86 1388.42 1063.78 1393.04 ;
     RECT  1074.14 1391.98 1117.06 1393.04 ;
     RECT  1173.98 1385.68 1210.18 1393.24 ;
     RECT  492.86 1393.04 1117.06 1394.16 ;
     RECT  349.34 1391.6 477.22 1399.58 ;
     RECT  349.82 1399.58 477.22 1400 ;
     RECT  1176.38 1393.24 1176.58 1400.8 ;
     RECT  349.82 1400 476.74 1405.04 ;
     RECT  293.18 1409.46 293.38 1409.88 ;
     RECT  494.78 1394.16 1117.06 1409.92 ;
     RECT  285.5 1409.88 293.38 1410.3 ;
     RECT  494.3 1409.92 1117.06 1412.86 ;
     RECT  285.02 1410.3 293.38 1414.08 ;
     RECT  349.82 1405.04 476.26 1417.86 ;
     RECT  285.02 1414.08 302.02 1418.28 ;
     RECT  349.34 1417.86 476.26 1418.48 ;
     RECT  285.02 1418.28 305.38 1418.9 ;
     RECT  -70 1349 219.46 1419 ;
     RECT  1588.185 1349 1870 1419 ;
     RECT  492.38 1412.86 1117.06 1422.52 ;
     RECT  301.82 1418.9 305.38 1422.9 ;
     RECT  349.34 1418.48 474.82 1424.58 ;
     RECT  488.54 1422.52 1117.06 1424.82 ;
     RECT  488.54 1424.82 877.54 1425.24 ;
     RECT  301.82 1422.9 307.3 1425.62 ;
     RECT  347.9 1424.58 474.82 1425.62 ;
     RECT  888.38 1424.82 1117.06 1425.7 ;
     RECT  347.9 1425.62 473.86 1426.68 ;
     RECT  1574.78 1385.68 1576.9 1426.84 ;
     RECT  285.02 1418.9 291.94 1429.2 ;
     RECT  301.82 1425.62 302.5 1429.2 ;
     RECT  346.94 1426.68 473.86 1429.62 ;
     RECT  0 1419 219.46 1437 ;
     RECT  1588.185 1419 1800 1437 ;
     RECT  285.02 1429.2 302.5 1437.38 ;
     RECT  291.26 1437.38 302.5 1439.7 ;
     RECT  313.34 1425.84 313.54 1439.7 ;
     RECT  291.26 1439.7 313.54 1440.54 ;
     RECT  341.18 1429.62 473.86 1440.54 ;
     RECT  291.26 1440.54 314.02 1440.96 ;
     RECT  341.18 1440.54 476.74 1444.52 ;
     RECT  273.5 1439.7 280.9 1444.74 ;
     RECT  341.18 1444.52 402.34 1445.16 ;
     RECT  291.26 1440.96 314.5 1445.58 ;
     RECT  340.7 1445.16 402.34 1445.58 ;
     RECT  270.14 1444.74 280.9 1447.26 ;
     RECT  291.26 1445.58 315.94 1447.26 ;
     RECT  333.02 1445.58 402.34 1447.26 ;
     RECT  413.18 1444.52 476.74 1447.46 ;
     RECT  488.54 1425.24 876.1 1447.5 ;
     RECT  263.9 1447.26 280.9 1447.68 ;
     RECT  413.18 1447.46 460.9 1447.88 ;
     RECT  255.74 1447.68 280.9 1448.1 ;
     RECT  291.26 1447.26 402.34 1448.1 ;
     RECT  413.18 1447.88 459.94 1448.3 ;
     RECT  456.38 1448.3 459.94 1452.08 ;
     RECT  255.74 1448.1 402.34 1454.82 ;
     RECT  255.74 1454.82 403.3 1456.92 ;
     RECT  413.18 1448.3 443.14 1456.92 ;
     RECT  476.54 1447.46 476.74 1457.72 ;
     RECT  490.94 1447.5 876.1 1458.42 ;
     RECT  460.22 1458.14 460.42 1458.56 ;
     RECT  471.26 1457.72 476.74 1458.56 ;
     RECT  255.74 1456.92 443.14 1459.86 ;
     RECT  233.66 1327.34 244.42 1460.44 ;
     RECT  490.94 1458.42 862.66 1461.36 ;
     RECT  490.94 1461.36 824.26 1462.2 ;
     RECT  837.5 1461.36 862.66 1462.62 ;
     RECT  846.62 1462.62 857.38 1463.04 ;
     RECT  501.5 1462.2 822.82 1463.46 ;
     RECT  490.94 1462.2 491.14 1465.14 ;
     RECT  846.62 1463.04 856.9 1465.56 ;
     RECT  501.5 1463.46 819.46 1465.98 ;
     RECT  846.62 1465.56 853.06 1465.98 ;
     RECT  254.78 1459.86 443.14 1466.36 ;
     RECT  501.5 1465.98 812.74 1466.4 ;
     RECT  846.62 1465.98 846.82 1466.4 ;
     RECT  254.78 1466.36 332.74 1467.62 ;
     RECT  347.42 1466.36 443.14 1467.84 ;
     RECT  260.06 1467.62 332.74 1468.04 ;
     RECT  501.5 1466.4 808.9 1468.92 ;
     RECT  502.46 1468.92 808.9 1469.34 ;
     RECT  502.46 1469.34 806.98 1470.18 ;
     RECT  260.06 1468.04 303.94 1470.56 ;
     RECT  318.14 1468.04 332.74 1470.56 ;
     RECT  721.82 1470.18 798.82 1470.6 ;
     RECT  260.06 1470.56 261.22 1470.98 ;
     RECT  273.5 1470.56 303.94 1470.98 ;
     RECT  318.62 1470.56 332.74 1470.98 ;
     RECT  502.46 1470.18 708.58 1471.02 ;
     RECT  283.58 1470.98 303.46 1471.4 ;
     RECT  324.86 1470.98 332.74 1471.4 ;
     RECT  460.22 1458.56 476.74 1471.4 ;
     RECT  721.82 1470.6 794.98 1471.44 ;
     RECT  260.06 1470.98 260.26 1471.82 ;
     RECT  273.5 1470.98 273.7 1471.82 ;
     RECT  347.42 1467.84 445.54 1471.82 ;
     RECT  347.42 1471.82 362.98 1472.24 ;
     RECT  708.38 1471.02 708.58 1472.28 ;
     RECT  502.46 1471.02 692.26 1472.7 ;
     RECT  721.82 1471.44 729.22 1472.7 ;
     RECT  834.62 1472.42 834.82 1472.84 ;
     RECT  691.58 1472.7 692.26 1473.12 ;
     RECT  745.82 1471.44 794.98 1473.12 ;
     RECT  502.46 1472.7 681.22 1473.54 ;
     RECT  721.82 1472.7 728.26 1473.54 ;
     RECT  745.82 1473.12 794.02 1473.54 ;
     RECT  324.86 1471.4 330.34 1473.92 ;
     RECT  502.94 1473.54 681.22 1473.96 ;
     RECT  721.82 1473.54 722.02 1473.96 ;
     RECT  745.82 1473.54 749.86 1473.96 ;
     RECT  760.7 1473.54 794.02 1473.96 ;
     RECT  347.42 1472.24 356.74 1474.34 ;
     RECT  764.06 1473.96 786.82 1474.38 ;
     RECT  285.02 1471.4 303.46 1475.18 ;
     RECT  347.42 1474.34 356.26 1475.18 ;
     RECT  372.86 1471.82 445.54 1475.18 ;
     RECT  692.06 1473.12 692.26 1475.22 ;
     RECT  286.94 1475.18 287.14 1475.6 ;
     RECT  299.9 1475.18 303.46 1475.6 ;
     RECT  433.34 1475.18 445.54 1475.82 ;
     RECT  324.86 1473.92 325.06 1476.02 ;
     RECT  627.26 1473.96 675.46 1476.48 ;
     RECT  528.86 1473.96 617.38 1477.32 ;
     RECT  627.26 1476.48 672.58 1477.32 ;
     RECT  764.06 1474.38 772.42 1477.32 ;
     RECT  502.94 1473.96 518.5 1477.74 ;
     RECT  561.5 1477.32 617.38 1477.74 ;
     RECT  627.26 1477.32 672.1 1477.74 ;
     RECT  770.3 1477.32 770.5 1477.74 ;
     RECT  433.34 1475.82 449.86 1478.12 ;
     RECT  502.94 1477.74 503.14 1478.16 ;
     RECT  636.86 1477.74 672.1 1478.16 ;
     RECT  378.62 1475.18 422.5 1478.54 ;
     RECT  433.34 1478.12 442.18 1478.54 ;
     RECT  528.86 1477.32 550.66 1478.58 ;
     RECT  414.14 1478.54 422.02 1478.96 ;
     RECT  433.82 1478.54 442.18 1478.96 ;
     RECT  381.98 1478.54 389.38 1479.38 ;
     RECT  402.62 1478.54 402.82 1479.38 ;
     RECT  414.14 1478.96 417.7 1479.38 ;
     RECT  433.82 1478.96 438.34 1479.38 ;
     RECT  -70 1437 219.46 1479.76 ;
     RECT  888.38 1425.7 1116.58 1480.18 ;
     RECT  528.86 1478.58 545.86 1480.26 ;
     RECT  569.66 1477.74 617.38 1480.26 ;
     RECT  573.98 1480.26 616.9 1480.68 ;
     RECT  666.14 1478.16 672.1 1480.68 ;
     RECT  518.3 1477.74 518.5 1481.1 ;
     RECT  528.86 1480.26 537.7 1481.1 ;
     RECT  577.34 1480.68 614.5 1481.1 ;
     RECT  636.86 1478.16 644.26 1481.1 ;
     RECT  666.14 1480.68 670.66 1481.1 ;
     RECT  528.86 1481.1 535.3 1481.52 ;
     RECT  577.82 1481.1 614.5 1481.52 ;
     RECT  666.14 1481.1 666.34 1481.52 ;
     RECT  528.86 1481.52 531.94 1481.94 ;
     RECT  580.7 1481.52 614.5 1481.94 ;
     RECT  636.86 1481.1 641.38 1481.94 ;
     RECT  529.82 1481.94 530.02 1482.36 ;
     RECT  580.7 1481.94 609.7 1482.36 ;
     RECT  580.7 1482.36 594.82 1482.66 ;
     RECT  580.7 1482.66 594.34 1484.88 ;
     RECT  581.66 1484.88 590.98 1485.3 ;
     RECT  590.78 1485.3 590.98 1485.72 ;
     RECT  233.66 1460.44 240.58 1493.84 ;
     RECT  273.02 1487.12 273.22 1493.84 ;
     RECT  1575.26 1426.84 1576.9 1497.7 ;
     RECT  -70 1479.76 211.815 1507 ;
     RECT  1588.185 1437 1870 1507 ;
     RECT  253.82 1486.7 254.02 1508.12 ;
     RECT  273.02 1493.84 280.42 1508.12 ;
     RECT  1575.26 1497.7 1576.42 1512.94 ;
     RECT  1575.26 1512.94 1575.46 1514.2 ;
     RECT  901.08 1480.18 1116.58 1524.28 ;
     RECT  0 1507 211.815 1525 ;
     RECT  1588.185 1507 1800 1525 ;
     RECT  901.08 1524.28 1085.38 1527.22 ;
     RECT  232.22 1493.84 240.58 1529.96 ;
     RECT  253.82 1508.12 280.42 1530.8 ;
     RECT  297.02 1494.26 297.22 1530.8 ;
     RECT  901.08 1527.22 1082.5 1535.2 ;
     RECT  253.82 1530.8 297.22 1537.52 ;
     RECT  971.9 1535.2 1082.5 1539.2 ;
     RECT  1098.62 1524.28 1116.58 1539.2 ;
     RECT  225.02 1529.96 240.58 1544.24 ;
     RECT  888.38 1480.18 890.02 1547.36 ;
     RECT  901.08 1535.2 961.54 1547.6 ;
     RECT  971.9 1539.2 1116.58 1547.6 ;
     RECT  901.08 1547.6 1116.58 1548.22 ;
     RECT  901.08 1548.22 1101.7 1549.48 ;
     RECT  901.08 1549.48 1083.94 1549.9 ;
     RECT  901.08 1549.9 1082.02 1554.52 ;
     RECT  1114.94 1548.22 1116.58 1554.94 ;
     RECT  918.14 1554.52 952.42 1560.82 ;
     RECT  918.62 1560.82 952.42 1561.66 ;
     RECT  924.38 1561.66 950.98 1562.08 ;
     RECT  927.26 1562.08 947.14 1562.5 ;
     RECT  927.26 1562.5 939.94 1569.64 ;
     RECT  966.62 1554.52 1082.02 1572.58 ;
     RECT  966.62 1572.58 1076.74 1573 ;
     RECT  966.62 1573 1074.34 1573.42 ;
     RECT  969.02 1573.42 1037.86 1575.94 ;
     RECT  969.98 1575.94 1037.86 1576.36 ;
     RECT  1047.74 1573.42 1074.34 1576.78 ;
     RECT  888.86 1547.36 890.02 1577.2 ;
     RECT  969.98 1576.36 1034.98 1577.2 ;
     RECT  1047.74 1576.78 1072.42 1577.2 ;
     RECT  253.82 1537.52 299.62 1577.42 ;
     RECT  889.82 1577.2 890.02 1577.62 ;
     RECT  981.98 1577.2 996.765 1577.62 ;
     RECT  222.62 1544.24 240.58 1577.88 ;
     RECT  251.42 1577.42 299.62 1577.88 ;
     RECT  320.06 1577 320.26 1577.88 ;
     RECT  1022.78 1577.2 1022.98 1578.04 ;
     RECT  222.62 1577.88 299.62 1578.1 ;
     RECT  320.06 1577.88 323.62 1578.1 ;
     RECT  222.62 1578.1 326.02 1578.26 ;
     RECT  222.62 1578.26 327.94 1578.46 ;
     RECT  1047.74 1577.2 1052.74 1578.46 ;
     RECT  222.62 1578.46 326.02 1578.82 ;
     RECT  261.02 1578.82 268.42 1579.3 ;
     RECT  268.22 1579.3 268.42 1579.72 ;
     RECT  311.235 1578.82 320.26 1579.72 ;
     RECT  786.62 1474.38 786.82 1579.895 ;
     RECT  901.08 1554.52 907.78 1579.895 ;
     RECT  -70 1525 211.815 1580.185 ;
     RECT  379.235 1579.895 384.765 1580.185 ;
     RECT  583.235 1579.895 588.765 1580.185 ;
     RECT  786.62 1579.895 792.765 1580.185 ;
     RECT  897.08 1579.895 907.78 1580.185 ;
     RECT  991.235 1577.62 996.765 1580.185 ;
     RECT  1186.46 1393.24 1210.18 1580.185 ;
     RECT  1399.235 1386.32 1405.54 1580.185 ;
     RECT  1588.185 1525 1870 1580.185 ;
     RECT  1012.7 1577.2 1012.9 1580.98 ;
     RECT  1051.58 1578.46 1052.74 1581.4 ;
     RECT  860.54 1580.78 860.74 1581.82 ;
     RECT  666.62 1558.52 666.82 1582.24 ;
     RECT  901.08 1580.185 907.78 1582.24 ;
     RECT  1051.58 1581.4 1051.78 1582.24 ;
     RECT  1116.38 1554.94 1116.58 1582.24 ;
     RECT  460.22 1471.4 471.46 1583.08 ;
     RECT  922.46 1577 922.66 1583.675 ;
     RECT  202.185 1580.185 211.815 1583.965 ;
     RECT  311.235 1579.72 316.765 1583.965 ;
     RECT  515.235 1583.675 520.765 1583.965 ;
     RECT  719.235 1583.675 724.765 1583.965 ;
     RECT  901.08 1582.24 902.92 1583.965 ;
     RECT  922.46 1583.675 928.765 1583.965 ;
     RECT  1127.235 1391.98 1140.1 1583.965 ;
     RECT  1331.235 1332.76 1336.765 1583.965 ;
     RECT  1535.235 1378.96 1540.765 1583.965 ;
     RECT  1588.185 1580.185 1597.815 1583.965 ;
     RECT  -70 1580.185 178 1595 ;
     RECT  1622 1580.185 1870 1595 ;
     RECT  922.46 1583.965 922.66 1598.3 ;
     RECT  922.46 1598.3 925.54 1598.5 ;
     RECT  749.66 1473.96 749.86 1601.78 ;
     RECT  925.34 1598.5 925.54 1616.06 ;
     RECT  1277.66 1361.54 1277.86 1616.06 ;
     RECT  414.14 1479.38 414.34 1619.42 ;
     RECT  0 1595 178 1620 ;
     RECT  414.14 1619.42 417.7 1620 ;
     RECT  506.3 1619.42 506.5 1620 ;
     RECT  593.18 1619.42 593.38 1620 ;
     RECT  677.66 1619.42 677.86 1620 ;
     RECT  748.7 1601.78 749.86 1620 ;
     RECT  786.62 1580.185 786.82 1620 ;
     RECT  834.62 1472.84 837.7 1620 ;
     RECT  875.9 1458.42 876.1 1620 ;
     RECT  924.86 1616.06 925.54 1620 ;
     RECT  1012.7 1603.04 1012.9 1620 ;
     RECT  1098.62 1549.48 1101.7 1620 ;
     RECT  1139.9 1583.965 1140.1 1620 ;
     RECT  1186.46 1580.185 1190.02 1620 ;
     RECT  1228.22 1393.04 1228.42 1620 ;
     RECT  1274.3 1616.06 1277.86 1620 ;
     RECT  1316.06 1392.62 1316.26 1620 ;
     RECT  1362.62 1363.22 1365.7 1620 ;
     RECT  1405.34 1580.185 1405.54 1620 ;
     RECT  1622 1595 1800 1620 ;
     RECT  1051.725 1620 1052.225 1620.045 ;
     RECT  0 1620 180 1622 ;
     RECT  414.14 1620 417.855 1622 ;
     RECT  502.145 1620 506.5 1622 ;
     RECT  590.145 1620 593.855 1622 ;
     RECT  677.66 1620 681.855 1622 ;
     RECT  746.225 1620 749.86 1622 ;
     RECT  786.62 1620 788.225 1622 ;
     RECT  834.225 1620 837.775 1622 ;
     RECT  875.725 1620 876.225 1622 ;
     RECT  922.225 1620 925.775 1622 ;
     RECT  963.725 1620 964.225 1622 ;
     RECT  1010.225 1620 1013.775 1622 ;
     RECT  1051.725 1620.045 1052.74 1622 ;
     RECT  1098.225 1620 1101.775 1622 ;
     RECT  1139.725 1620 1140.225 1622 ;
     RECT  1186.225 1620 1190.02 1622 ;
     RECT  1209.98 1580.185 1210.18 1622 ;
     RECT  1227.725 1620 1228.42 1622 ;
     RECT  1274.225 1620 1277.86 1622 ;
     RECT  1315.725 1620 1316.26 1622 ;
     RECT  1362.225 1620 1365.775 1622 ;
     RECT  1403.725 1620 1405.54 1622 ;
     RECT  1620 1620 1800 1622 ;
     RECT  0 1622 1800 1800 ;
     RECT  205 1800 275 1870 ;
     RECT  293 1800 363 1870 ;
     RECT  381 1800 451 1870 ;
     RECT  469 1800 539 1870 ;
     RECT  557 1800 627 1870 ;
     RECT  645 1800 715 1870 ;
     RECT  733 1800 803 1870 ;
     RECT  821 1800 891 1870 ;
     RECT  909 1800 979 1870 ;
     RECT  997 1800 1067 1870 ;
     RECT  1085 1800 1155 1870 ;
     RECT  1173 1800 1243 1870 ;
     RECT  1261 1800 1331 1870 ;
     RECT  1349 1800 1419 1870 ;
     RECT  1437 1800 1507 1870 ;
     RECT  1525 1800 1595 1870 ;
    LAYER Metal4 ;
     RECT  -70 205 0 275 ;
     RECT  -70 293 0 363 ;
     RECT  -70 381 0 451 ;
     RECT  -70 469 0 539 ;
     RECT  -70 557 0 627 ;
     RECT  -70 645 0 715 ;
     RECT  -70 733 0 803 ;
     RECT  -70 821 0 891 ;
     RECT  -70 909 0 979 ;
     RECT  -70 997 0 1067 ;
     RECT  -70 1085 0 1155 ;
     RECT  -70 1173 0 1243 ;
     RECT  -70 1261 0 1331 ;
     RECT  -70 1349 0 1419 ;
     RECT  -70 1437 0 1507 ;
     RECT  -70 1525 0 1595 ;
     RECT  0 0 178 1800 ;
     RECT  178 0 180 180 ;
     RECT  178 1620 180 1800 ;
     RECT  178 219.14 202.14 1580.14 ;
     RECT  180 0 205 178 ;
     RECT  180 1622 205 1800 ;
     RECT  202.14 215.36 211.86 1583.92 ;
     RECT  211.86 422.15 233.66 551.33 ;
     RECT  211.86 944.06 233.86 944.26 ;
     RECT  229.34 647.54 235.1 647.74 ;
     RECT  233.66 422.15 236.26 552.4 ;
     RECT  236.06 1449.32 236.54 1449.52 ;
     RECT  211.86 613.94 237.02 614.14 ;
     RECT  237.02 613.94 239.9 619.18 ;
     RECT  224.06 634.52 239.9 634.72 ;
     RECT  211.86 1207.82 240.58 1208.02 ;
     RECT  235.58 383.36 241.34 383.56 ;
     RECT  211.86 1301.06 241.34 1301.26 ;
     RECT  211.86 855.86 241.82 856.06 ;
     RECT  235.58 1343.06 241.82 1343.26 ;
     RECT  211.86 704.05 242.3 833.23 ;
     RECT  241.82 855.86 242.3 866.56 ;
     RECT  241.82 1335.08 242.3 1343.26 ;
     RECT  242.3 855.86 242.78 866.98 ;
     RECT  242.3 1335.08 242.78 1344.94 ;
     RECT  242.3 702.98 243.26 833.23 ;
     RECT  236.54 1449.32 243.26 1449.94 ;
     RECT  243.26 1449.32 243.74 1458.34 ;
     RECT  242.78 852.92 244.22 866.98 ;
     RECT  243.74 1449.32 244.22 1460.02 ;
     RECT  237.02 1468.64 244.22 1468.84 ;
     RECT  244.7 1220.42 246.82 1220.62 ;
     RECT  243.26 702.98 247.58 838.84 ;
     RECT  243.74 656.78 248.06 656.98 ;
     RECT  248.06 1051.62 248.54 1051.82 ;
     RECT  245.66 1172.58 248.54 1172.78 ;
     RECT  244.22 852.92 249.02 867.82 ;
     RECT  236.26 422.15 249.98 551.33 ;
     RECT  249.98 1110.42 250.46 1110.62 ;
     RECT  245.18 1119.62 250.46 1119.82 ;
     RECT  250.46 1110.42 250.66 1119.82 ;
     RECT  248.54 1169.22 251.42 1172.78 ;
     RECT  240.38 1574.06 251.42 1574.26 ;
     RECT  250.66 1110.42 251.62 1113.98 ;
     RECT  249.98 420.74 252.38 551.33 ;
     RECT  251.42 1168.8 252.86 1172.78 ;
     RECT  252.38 419.06 253.34 551.33 ;
     RECT  248.54 1047.42 253.34 1051.82 ;
     RECT  252.86 1168.8 253.34 1176.14 ;
     RECT  240.86 1285.1 253.34 1285.3 ;
     RECT  253.34 1047.42 253.54 1052.66 ;
     RECT  253.34 1168.8 253.82 1182.44 ;
     RECT  253.34 1285.1 254.02 1286.6 ;
     RECT  211.86 1031 254.78 1031.2 ;
     RECT  254.3 1224.66 254.78 1224.86 ;
     RECT  251.42 1089.84 254.98 1090.04 ;
     RECT  243.74 878.12 255.26 878.32 ;
     RECT  250.94 1065.44 255.46 1065.64 ;
     RECT  253.34 419.06 255.94 551.98 ;
     RECT  253.82 1161.24 255.94 1182.44 ;
     RECT  254.78 1224.66 255.94 1226.12 ;
     RECT  234.62 1515.26 256.22 1515.46 ;
     RECT  255.94 1224.66 256.42 1225.7 ;
     RECT  241.34 1301.06 256.7 1306.72 ;
     RECT  253.82 1191.06 256.9 1191.26 ;
     RECT  253.54 1048.26 257.18 1052.66 ;
     RECT  255.94 1168.8 257.18 1182.44 ;
     RECT  251.62 1113.78 257.38 1113.98 ;
     RECT  256.42 1225.5 257.38 1225.7 ;
     RECT  255.94 419.06 258.14 551.33 ;
     RECT  251.42 1574.06 258.14 1577.62 ;
     RECT  249.02 852.92 258.62 868.24 ;
     RECT  255.26 877.28 258.62 878.32 ;
     RECT  258.14 1574.06 258.62 1582.66 ;
     RECT  258.14 1203.66 259.58 1203.86 ;
     RECT  256.7 1301.06 259.58 1312.64 ;
     RECT  250.94 1099.5 260.06 1099.7 ;
     RECT  257.18 1168.8 262.18 1187.48 ;
     RECT  254.02 1285.1 262.46 1285.3 ;
     RECT  254.78 1026 262.66 1031.2 ;
     RECT  257.18 1048.26 262.66 1053.92 ;
     RECT  260.06 1098.24 262.66 1099.7 ;
     RECT  262.46 1123.02 262.94 1123.22 ;
     RECT  259.58 1296.9 263.42 1312.64 ;
     RECT  256.22 1508.54 263.42 1515.46 ;
     RECT  260.06 1010.04 263.9 1010.24 ;
     RECT  262.94 1100.76 263.9 1100.96 ;
     RECT  257.66 675.68 264.38 675.88 ;
     RECT  263.9 1100.76 264.38 1101.8 ;
     RECT  263.9 1110.42 264.38 1110.62 ;
     RECT  254.78 689.12 264.86 689.32 ;
     RECT  247.58 701.3 264.86 838.84 ;
     RECT  262.94 1123.02 264.86 1127.42 ;
     RECT  256.22 1137.72 264.86 1137.92 ;
     RECT  262.46 1278 265.06 1285.3 ;
     RECT  263.42 1293.96 265.06 1315.58 ;
     RECT  262.66 1048.26 265.34 1048.46 ;
     RECT  261.98 1078.08 265.34 1078.28 ;
     RECT  262.18 1172.58 265.34 1187.48 ;
     RECT  259.58 1196.52 265.34 1203.86 ;
     RECT  264.86 1123.02 265.54 1137.92 ;
     RECT  263.42 1508.12 265.82 1515.46 ;
     RECT  265.34 1040.28 266.02 1048.46 ;
     RECT  265.34 1172.58 266.5 1203.86 ;
     RECT  265.06 1293.96 266.5 1314.74 ;
     RECT  264.38 1100.76 266.98 1110.62 ;
     RECT  265.34 1074.3 267.26 1078.28 ;
     RECT  263.9 1009.2 267.94 1010.24 ;
     RECT  266.78 1039.02 267.94 1039.22 ;
     RECT  258.14 418.64 269.18 551.33 ;
     RECT  267.26 1074.3 269.38 1082.06 ;
     RECT  266.98 1100.76 269.38 1107.68 ;
     RECT  266.5 1293.96 269.38 1312.64 ;
     RECT  268.22 1153.68 269.86 1153.88 ;
     RECT  267.74 1240.62 270.14 1240.82 ;
     RECT  266.78 992.4 270.34 992.6 ;
     RECT  267.94 1010.04 270.34 1010.24 ;
     RECT  262.66 1026 270.34 1026.2 ;
     RECT  266.02 1048.26 270.34 1048.46 ;
     RECT  267.74 1059.6 270.62 1059.8 ;
     RECT  270.14 1068.84 270.62 1069.04 ;
     RECT  269.38 1081.44 270.62 1082.06 ;
     RECT  270.14 1209.96 270.62 1210.16 ;
     RECT  258.62 1574.06 270.62 1583.08 ;
     RECT  270.62 1081.44 271.1 1089.62 ;
     RECT  270.62 1059.6 271.3 1069.04 ;
     RECT  271.1 1081.44 271.3 1100.54 ;
     RECT  265.54 1123.02 271.3 1130.78 ;
     RECT  270.14 1240.62 271.3 1241.66 ;
     RECT  248.06 656.78 271.58 663.28 ;
     RECT  271.3 1059.6 271.58 1066.94 ;
     RECT  271.3 1123.02 271.58 1123.22 ;
     RECT  270.62 1209.96 271.58 1215.2 ;
     RECT  271.3 1081.44 271.78 1082.06 ;
     RECT  271.58 1122.18 271.78 1123.22 ;
     RECT  269.38 1297.74 271.78 1312.64 ;
     RECT  239.9 613.94 272.06 634.72 ;
     RECT  266.5 1172.58 272.06 1197.98 ;
     RECT  272.06 1169.64 272.26 1197.98 ;
     RECT  271.78 1297.74 272.26 1308.86 ;
     RECT  235.1 647.12 272.54 647.74 ;
     RECT  271.58 656.78 272.54 666.22 ;
     RECT  242.78 1335.08 272.54 1345.78 ;
     RECT  272.26 1189.38 272.74 1197.98 ;
     RECT  253.82 1486.7 273.02 1486.9 ;
     RECT  271.78 1081.44 273.22 1081.64 ;
     RECT  272.26 1298.58 273.22 1308.86 ;
     RECT  271.58 1209.96 274.46 1221.08 ;
     RECT  274.46 1209.96 274.94 1221.5 ;
     RECT  265.06 1278.42 274.94 1285.3 ;
     RECT  205 -70 275 178 ;
     RECT  205 1622 275 1870 ;
     RECT  273.02 1236.84 275.14 1237.04 ;
     RECT  274.46 976.02 275.42 976.22 ;
     RECT  270.14 1152.84 275.42 1153.04 ;
     RECT  272.74 1191.9 275.42 1197.98 ;
     RECT  274.94 1206.6 275.42 1221.5 ;
     RECT  253.82 1255.32 275.42 1255.52 ;
     RECT  225.02 1529.96 275.42 1530.16 ;
     RECT  271.3 1093.62 275.62 1100.54 ;
     RECT  274.94 1271.28 275.62 1285.3 ;
     RECT  275.62 1100.34 276.1 1100.54 ;
     RECT  275.42 976.02 277.06 980.42 ;
     RECT  273.22 1298.58 277.54 1306.72 ;
     RECT  272.54 1327.14 277.54 1345.78 ;
     RECT  265.82 1508.12 277.82 1515.88 ;
     RECT  277.54 1333.82 278.02 1345.78 ;
     RECT  277.82 1107.9 278.3 1108.1 ;
     RECT  276.38 1021.38 278.5 1021.58 ;
     RECT  272.26 1169.64 278.78 1180.34 ;
     RECT  275.42 1255.32 278.78 1259.3 ;
     RECT  278.78 1168.8 279.46 1180.34 ;
     RECT  275.42 1191.9 279.94 1221.5 ;
     RECT  273.02 1486.7 280.22 1487.32 ;
     RECT  277.82 1500.98 280.22 1515.88 ;
     RECT  277.06 978.96 280.42 980.42 ;
     RECT  269.18 418.22 280.7 551.33 ;
     RECT  271.78 1122.18 281.18 1122.38 ;
     RECT  278.78 1255.32 281.18 1260.56 ;
     RECT  275.62 1271.28 281.18 1271.48 ;
     RECT  279.94 1191.9 281.38 1221.08 ;
     RECT  278.3 1107.9 282.14 1112.3 ;
     RECT  281.18 1122.18 282.14 1130.78 ;
     RECT  280.42 979.38 282.34 980.42 ;
     RECT  277.82 1031.46 282.82 1031.66 ;
     RECT  271.58 1051.2 282.82 1066.94 ;
     RECT  281.38 1206.6 282.82 1221.08 ;
     RECT  282.14 1233.9 283.3 1234.1 ;
     RECT  283.1 1073.46 283.58 1073.66 ;
     RECT  275.42 1150.74 283.58 1153.04 ;
     RECT  279.46 1168.8 283.78 1169 ;
     RECT  281.38 1191.9 284.26 1195.88 ;
     RECT  282.62 1551.38 285.02 1551.58 ;
     RECT  282.14 1107.9 285.98 1130.78 ;
     RECT  279.46 1178.46 286.46 1180.34 ;
     RECT  284.26 1191.9 286.46 1192.1 ;
     RECT  281.18 1255.32 286.94 1271.48 ;
     RECT  275.62 1285.1 286.94 1285.3 ;
     RECT  272.54 647.12 287.42 666.22 ;
     RECT  282.82 1051.2 287.62 1061.06 ;
     RECT  264.86 689.12 287.9 838.84 ;
     RECT  277.54 1299.42 287.9 1306.72 ;
     RECT  285.98 1319.58 287.9 1319.78 ;
     RECT  286.94 986.94 288.1 987.14 ;
     RECT  283.58 1150.74 288.38 1158.08 ;
     RECT  287.62 1053.3 288.58 1061.06 ;
     RECT  286.94 1255.32 288.58 1285.3 ;
     RECT  284.54 1031.88 288.86 1032.08 ;
     RECT  288.86 1031.88 289.06 1037.54 ;
     RECT  288.58 1053.3 289.06 1060.64 ;
     RECT  288.38 1142.34 289.06 1165.22 ;
     RECT  275.42 1529.96 289.82 1530.58 ;
     RECT  289.06 1053.3 290.02 1060.22 ;
     RECT  289.06 1150.32 290.02 1165.22 ;
     RECT  285.98 1106.22 290.3 1130.78 ;
     RECT  282.82 1206.6 290.78 1219.4 ;
     RECT  264.38 675.68 291.26 676.3 ;
     RECT  287.9 687.86 291.26 838.84 ;
     RECT  288.38 1005.84 291.74 1006.04 ;
     RECT  290.3 1106.22 292.22 1138.34 ;
     RECT  289.82 1529.96 292.22 1531 ;
     RECT  285.02 1544.24 292.22 1551.58 ;
     RECT  286.46 1178.46 292.7 1192.1 ;
     RECT  275 0 293 178 ;
     RECT  275 1622 293 1800 ;
     RECT  292.22 1104.54 293.18 1138.34 ;
     RECT  290.78 1206.18 293.66 1219.4 ;
     RECT  278.02 1333.82 293.66 1334.48 ;
     RECT  278.02 1343.06 293.66 1345.78 ;
     RECT  291.74 1002.06 293.86 1006.04 ;
     RECT  283.58 1073.46 294.14 1074.08 ;
     RECT  292.7 1176.36 295.1 1195.46 ;
     RECT  294.14 1073.46 295.3 1082.48 ;
     RECT  290.02 1150.32 295.3 1158.08 ;
     RECT  288.58 1271.28 295.3 1285.3 ;
     RECT  294.14 1238.94 295.78 1239.14 ;
     RECT  293.66 1333.82 296.74 1345.78 ;
     RECT  280.7 411.08 297.02 551.33 ;
     RECT  287.42 646.7 297.02 666.22 ;
     RECT  290.02 1053.3 297.22 1057.7 ;
     RECT  296.74 1333.82 297.22 1334.48 ;
     RECT  297.22 1053.3 297.7 1055.6 ;
     RECT  293.18 1100.34 297.7 1138.34 ;
     RECT  297.7 1100.34 298.94 1131.62 ;
     RECT  295.3 1150.74 298.94 1158.08 ;
     RECT  295.1 1167.96 298.94 1195.46 ;
     RECT  295.3 1276.74 298.94 1285.3 ;
     RECT  297.7 1055.4 299.14 1055.6 ;
     RECT  288.58 1255.32 299.42 1258.88 ;
     RECT  298.94 1096.98 299.62 1131.62 ;
     RECT  272.06 608.06 300.38 634.72 ;
     RECT  297.02 645.44 300.38 666.22 ;
     RECT  293.66 1206.18 301.34 1220.66 ;
     RECT  298.94 1276.74 301.34 1289.54 ;
     RECT  287.9 1299.42 301.34 1319.78 ;
     RECT  301.34 1206.18 301.54 1221.5 ;
     RECT  301.54 1207.44 301.82 1221.5 ;
     RECT  301.34 1276.74 302.02 1319.78 ;
     RECT  289.06 1037.34 302.3 1037.54 ;
     RECT  299.62 1096.98 302.3 1112.72 ;
     RECT  299.42 1250.28 302.78 1264.34 ;
     RECT  297.5 1233.06 302.98 1233.26 ;
     RECT  302.3 1091.94 303.46 1112.72 ;
     RECT  302.78 1243.98 303.46 1264.34 ;
     RECT  302.02 1276.74 303.46 1299.62 ;
     RECT  293.18 561.02 303.74 561.22 ;
     RECT  211.86 570.26 303.74 575.5 ;
     RECT  303.46 1243.98 304.42 1262.66 ;
     RECT  296.74 1343.06 304.42 1345.78 ;
     RECT  298.94 1150.74 305.18 1195.46 ;
     RECT  303.46 1276.74 305.38 1289.54 ;
     RECT  302.3 1036.92 305.66 1037.54 ;
     RECT  303.46 1107.9 306.34 1112.72 ;
     RECT  302.02 1312.02 306.34 1319.78 ;
     RECT  295.3 1073.46 306.62 1074.08 ;
     RECT  303.46 1091.94 306.82 1097.18 ;
     RECT  304.42 1343.06 306.82 1345.36 ;
     RECT  300.38 608.06 307.58 666.22 ;
     RECT  291.26 675.68 307.58 838.84 ;
     RECT  299.62 1122.18 308.06 1131.62 ;
     RECT  301.82 1207.44 308.06 1222.34 ;
     RECT  306.62 1073.46 308.26 1074.92 ;
     RECT  297.22 1333.82 308.26 1334.02 ;
     RECT  305.38 1276.74 308.74 1282.4 ;
     RECT  308.26 1073.46 309.22 1073.66 ;
     RECT  297.02 411.08 309.5 552.4 ;
     RECT  303.74 561.02 309.5 575.5 ;
     RECT  308.06 1121.34 309.5 1131.62 ;
     RECT  305.18 1145.7 309.5 1195.46 ;
     RECT  309.5 1121.34 309.7 1195.46 ;
     RECT  308.74 1276.74 309.7 1281.98 ;
     RECT  309.7 1281.36 310.66 1281.98 ;
     RECT  309.7 1122.18 311.14 1195.46 ;
     RECT  241.34 383.36 311.19 388.18 ;
     RECT  309.5 411.08 311.19 575.5 ;
     RECT  211.86 592.1 311.19 592.3 ;
     RECT  307.58 608.06 311.19 838.84 ;
     RECT  258.62 852.92 311.19 878.32 ;
     RECT  270.62 1573.22 311.19 1583.08 ;
     RECT  306.82 1343.06 311.62 1344.94 ;
     RECT  293.86 1005.84 311.9 1006.04 ;
     RECT  308.06 1207.44 312.1 1225.7 ;
     RECT  306.34 1111.68 313.34 1112.72 ;
     RECT  311.14 1184.76 313.54 1195.46 ;
     RECT  312.1 1207.86 313.54 1225.7 ;
     RECT  311.14 1139.82 314.02 1150.94 ;
     RECT  313.54 1217.94 314.02 1225.7 ;
     RECT  304.42 1243.98 314.02 1260.98 ;
     RECT  311.62 1343.06 314.02 1344.52 ;
     RECT  311.9 1005.84 314.78 1010.24 ;
     RECT  314.02 1243.98 314.78 1251.74 ;
     RECT  311.14 1122.18 314.98 1131.2 ;
     RECT  312.38 1327.56 314.98 1327.76 ;
     RECT  313.34 1111.68 315.26 1113.56 ;
     RECT  314.02 1139.82 315.94 1145.9 ;
     RECT  313.54 1191.48 315.94 1195.46 ;
     RECT  314.02 1343.06 316.42 1344.1 ;
     RECT  312.86 979.38 316.7 979.58 ;
     RECT  311.19 215.36 316.81 878.32 ;
     RECT  311.19 1573.22 316.81 1583.92 ;
     RECT  315.94 1193.16 316.9 1195.46 ;
     RECT  314.02 1217.94 316.9 1218.56 ;
     RECT  315.94 1139.82 317.38 1140.02 ;
     RECT  310.66 1281.36 317.38 1281.56 ;
     RECT  316.9 1217.94 317.86 1218.14 ;
     RECT  298.94 1429.2 317.86 1429.4 ;
     RECT  315.26 1104.12 318.14 1113.56 ;
     RECT  311.14 1165.44 318.34 1176.14 ;
     RECT  314.78 1002.06 318.62 1010.24 ;
     RECT  314.78 1235.58 318.82 1251.74 ;
     RECT  316.42 1343.48 318.82 1344.1 ;
     RECT  318.14 1104.12 319.3 1119.02 ;
     RECT  318.82 1235.58 320.54 1251.32 ;
     RECT  316.7 976.86 320.74 979.58 ;
     RECT  314.02 1260.36 320.74 1260.98 ;
     RECT  306.34 1312.02 320.74 1315.58 ;
     RECT  314.98 1130.58 321.22 1131.2 ;
     RECT  321.02 1054.98 321.98 1055.18 ;
     RECT  318.34 1165.44 321.98 1165.64 ;
     RECT  306.82 1091.94 323.42 1092.14 ;
     RECT  319.3 1104.12 323.42 1116.5 ;
     RECT  318.82 1343.9 323.62 1344.1 ;
     RECT  321.98 1157.88 324.1 1165.64 ;
     RECT  321.98 1054.98 324.38 1058.54 ;
     RECT  305.66 1036.92 325.34 1039.64 ;
     RECT  323.42 1091.94 326.02 1116.5 ;
     RECT  318.62 1002.06 326.3 1010.66 ;
     RECT  315.26 1024.74 326.3 1028.3 ;
     RECT  326.3 1002.06 326.78 1028.3 ;
     RECT  325.34 1036.92 326.78 1043 ;
     RECT  324.38 1052.04 326.78 1058.54 ;
     RECT  320.74 976.86 327.26 978.32 ;
     RECT  326.78 1002.06 327.26 1059.8 ;
     RECT  317.18 1074.3 327.26 1074.5 ;
     RECT  266.3 1359.06 327.26 1359.26 ;
     RECT  326.02 1104.96 327.46 1116.5 ;
     RECT  326.02 1091.94 327.74 1092.14 ;
     RECT  320.54 1230.54 327.74 1251.32 ;
     RECT  320.74 1260.36 327.74 1260.56 ;
     RECT  327.26 1002.06 328.7 1074.5 ;
     RECT  327.26 968.46 329.18 978.32 ;
     RECT  313.54 1207.86 329.18 1208.06 ;
     RECT  327.74 1230.54 329.18 1260.56 ;
     RECT  329.18 963.42 329.66 978.32 ;
     RECT  316.9 1193.16 329.66 1193.36 ;
     RECT  327.46 1104.96 330.34 1110.2 ;
     RECT  329.18 1229.28 330.34 1260.56 ;
     RECT  328.22 1147.8 331.1 1148 ;
     RECT  329.18 1206.18 331.1 1208.06 ;
     RECT  316.81 411.08 331.58 551.33 ;
     RECT  330.34 1230.54 331.58 1260.56 ;
     RECT  320.54 1289.76 331.58 1289.96 ;
     RECT  303.46 1299.42 331.58 1299.62 ;
     RECT  322.46 1136.04 332.54 1136.24 ;
     RECT  331.1 1146.12 332.54 1148 ;
     RECT  329.66 960.9 332.74 978.32 ;
     RECT  332.54 1136.04 332.74 1148 ;
     RECT  332.74 1136.04 333.22 1138.34 ;
     RECT  332.74 1147.8 333.5 1148 ;
     RECT  324.1 1157.88 333.5 1159.76 ;
     RECT  331.58 1230.54 333.5 1261.82 ;
     RECT  332.74 963.42 333.7 978.32 ;
     RECT  333.5 1147.8 333.7 1159.76 ;
     RECT  333.22 1136.04 333.98 1136.24 ;
     RECT  329.66 1189.8 333.98 1193.36 ;
     RECT  331.1 1206.18 333.98 1210.58 ;
     RECT  328.7 1002.06 334.66 1081.22 ;
     RECT  328.22 990.72 334.94 990.92 ;
     RECT  333.7 968.46 335.14 978.32 ;
     RECT  316.81 592.1 335.42 592.3 ;
     RECT  331.58 1289.76 335.42 1299.62 ;
     RECT  335.42 1289.34 336.38 1299.62 ;
     RECT  330.34 1104.96 336.86 1109.78 ;
     RECT  333.98 1189.8 336.86 1210.58 ;
     RECT  336.38 1288.92 337.34 1299.62 ;
     RECT  334.66 1002.9 337.82 1081.22 ;
     RECT  327.74 1091.52 337.82 1092.14 ;
     RECT  336.86 1104.12 337.82 1109.78 ;
     RECT  334.94 1331.76 337.82 1331.96 ;
     RECT  333.5 1230.54 338.3 1263.08 ;
     RECT  326.78 1278 338.3 1278.2 ;
     RECT  337.34 1288.92 338.3 1300.88 ;
     RECT  336.86 1189.8 339.46 1217.3 ;
     RECT  337.82 1002.9 339.74 1109.78 ;
     RECT  339.74 1002.9 341.86 1110.62 ;
     RECT  337.82 1327.14 341.86 1331.96 ;
     RECT  341.86 1103.28 342.14 1110.62 ;
     RECT  340.7 1123.86 342.62 1124.06 ;
     RECT  333.98 1134.78 342.62 1136.24 ;
     RECT  338.3 1230.54 342.62 1300.88 ;
     RECT  341.66 931.08 342.82 931.28 ;
     RECT  335.14 978.12 342.82 978.32 ;
     RECT  337.34 1178.46 343.1 1178.66 ;
     RECT  342.62 1230.54 343.1 1306.76 ;
     RECT  342.14 1103.28 343.58 1111.04 ;
     RECT  341.86 1002.9 343.78 1092.14 ;
     RECT  335.14 968.46 344.06 968.66 ;
     RECT  334.94 990.72 344.06 994.28 ;
     RECT  343.1 1175.94 344.06 1178.66 ;
     RECT  331.58 411.08 344.54 551.98 ;
     RECT  316.81 560.6 344.54 575.5 ;
     RECT  333.7 1151.58 344.54 1159.76 ;
     RECT  344.06 1172.16 344.54 1178.66 ;
     RECT  343.1 1230.54 345.22 1312.22 ;
     RECT  342.62 1123.86 346.18 1136.24 ;
     RECT  345.22 1247.76 346.18 1271.06 ;
     RECT  344.54 1151.58 346.94 1178.66 ;
     RECT  339.46 1189.8 346.94 1210.58 ;
     RECT  344.06 965.52 347.14 968.66 ;
     RECT  346.18 1270.86 348.1 1271.06 ;
     RECT  343.58 1103.28 348.86 1114.4 ;
     RECT  346.18 1123.86 348.86 1131.62 ;
     RECT  345.22 1230.54 348.86 1236.2 ;
     RECT  211.86 1386.32 349.06 1386.52 ;
     RECT  346.94 1151.58 349.54 1210.58 ;
     RECT  343.78 1006.26 350.3 1092.14 ;
     RECT  348.86 1103.28 350.3 1131.62 ;
     RECT  349.54 1175.1 350.3 1210.58 ;
     RECT  345.22 1280.94 350.98 1312.22 ;
     RECT  344.54 411.08 351.26 575.5 ;
     RECT  350.98 1291.44 351.46 1312.22 ;
     RECT  348.86 1225.92 351.74 1236.2 ;
     RECT  351.74 1225.5 352.9 1236.2 ;
     RECT  347.14 968.46 353.18 968.66 ;
     RECT  350.3 1175.1 353.18 1211 ;
     RECT  349.34 926.88 353.38 927.08 ;
     RECT  344.06 990.72 353.38 994.7 ;
     RECT  341.86 1327.14 353.38 1331.54 ;
     RECT  353.18 1175.1 353.66 1211.42 ;
     RECT  353.18 968.46 353.86 969.5 ;
     RECT  353.66 1175.1 353.86 1213.1 ;
     RECT  350.98 1280.94 353.86 1281.98 ;
     RECT  350.3 1006.26 354.34 1131.62 ;
     RECT  352.9 1225.92 354.62 1236.2 ;
     RECT  346.94 1140.24 355.1 1140.86 ;
     RECT  349.54 1151.58 355.1 1165.22 ;
     RECT  353.38 1327.14 356.26 1330.7 ;
     RECT  355.58 1383 356.26 1383.2 ;
     RECT  353.86 1175.1 356.74 1212.26 ;
     RECT  346.18 1247.76 356.74 1262.24 ;
     RECT  354.62 1271.28 356.74 1271.48 ;
     RECT  351.46 1299.42 356.74 1312.22 ;
     RECT  316.81 383.36 357.02 388.18 ;
     RECT  356.74 1247.76 357.22 1261.82 ;
     RECT  357.22 1261.62 357.7 1261.82 ;
     RECT  357.02 383.36 357.98 389.02 ;
     RECT  354.34 1103.28 357.98 1131.62 ;
     RECT  355.1 1140.24 357.98 1165.22 ;
     RECT  327.26 1353.6 358.18 1359.26 ;
     RECT  357.98 383.36 358.46 395.32 ;
     RECT  356.54 949.14 358.46 949.34 ;
     RECT  353.86 1281.78 359.62 1281.98 ;
     RECT  357.22 1247.76 360.1 1251.32 ;
     RECT  356.54 926.46 360.38 926.66 ;
     RECT  358.46 949.14 361.06 950.18 ;
     RECT  360.38 984.84 361.34 985.04 ;
     RECT  354.62 1225.92 362.3 1237.04 ;
     RECT  361.34 983.58 362.78 985.04 ;
     RECT  353.38 994.5 362.78 994.7 ;
     RECT  356.26 1327.56 362.98 1330.7 ;
     RECT  293 -70 363 178 ;
     RECT  293 1622 363 1870 ;
     RECT  357.98 1103.28 363.26 1165.22 ;
     RECT  354.34 1006.26 363.74 1092.14 ;
     RECT  363.26 1103.28 363.74 1165.64 ;
     RECT  362.3 1221.3 363.74 1237.04 ;
     RECT  358.46 382.94 364.22 395.32 ;
     RECT  358.18 1359.06 364.22 1359.26 ;
     RECT  360.38 922.26 364.7 926.66 ;
     RECT  361.06 949.98 365.86 950.18 ;
     RECT  363.74 1221.3 366.62 1244.18 ;
     RECT  364.7 922.26 366.82 931.28 ;
     RECT  364.22 1359.06 367.3 1361.78 ;
     RECT  366.82 923.1 367.78 931.28 ;
     RECT  356.74 1175.1 368.06 1211 ;
     RECT  366.62 1220.88 368.06 1244.18 ;
     RECT  356.74 1312.02 368.06 1312.22 ;
     RECT  368.54 1289.76 369.02 1289.96 ;
     RECT  356.74 1299.42 369.02 1299.62 ;
     RECT  362.78 983.58 370.18 994.7 ;
     RECT  368.06 1175.1 370.46 1244.18 ;
     RECT  362.98 1330.5 370.66 1330.7 ;
     RECT  370.18 991.98 370.94 994.7 ;
     RECT  363.74 1006.26 370.94 1165.64 ;
     RECT  369.02 1289.76 370.94 1299.62 ;
     RECT  368.06 1309.08 370.94 1312.22 ;
     RECT  370.46 969.3 371.42 969.5 ;
     RECT  370.94 991.98 371.42 1165.64 ;
     RECT  370.46 1175.1 371.42 1244.6 ;
     RECT  370.94 1289.76 371.42 1314.74 ;
     RECT  371.42 1288.08 371.62 1314.74 ;
     RECT  371.42 991.98 372.1 1244.6 ;
     RECT  371.42 969.3 372.58 980.84 ;
     RECT  371.9 1411.14 372.58 1411.34 ;
     RECT  370.46 1273.38 372.86 1273.58 ;
     RECT  371.9 1331.34 372.86 1334.9 ;
     RECT  372.1 1006.26 373.34 1244.6 ;
     RECT  372.86 1255.32 373.34 1255.52 ;
     RECT  370.94 1381.74 373.34 1381.94 ;
     RECT  372.58 978.54 373.54 980.84 ;
     RECT  371.62 1288.08 374.02 1312.22 ;
     RECT  316.81 852.92 374.3 878.32 ;
     RECT  372.86 1272.96 374.3 1273.58 ;
     RECT  373.34 1380.06 374.3 1381.94 ;
     RECT  374.02 1289.76 374.98 1312.22 ;
     RECT  316.81 608.06 375.26 838.84 ;
     RECT  374.3 1380.06 375.26 1389.08 ;
     RECT  364.22 381.26 376.22 395.32 ;
     RECT  351.26 404.78 376.22 575.5 ;
     RECT  373.34 1006.26 376.42 1255.52 ;
     RECT  367.3 1359.06 376.7 1361.36 ;
     RECT  375.26 1376.28 376.7 1389.08 ;
     RECT  375.74 910.5 377.86 910.7 ;
     RECT  376.7 1359.06 378.62 1363.04 ;
     RECT  378.14 942.42 379.1 942.62 ;
     RECT  376.22 381.26 379.19 575.5 ;
     RECT  335.42 587.06 379.19 592.3 ;
     RECT  375.26 608.06 379.19 842.62 ;
     RECT  374.3 852.92 379.19 884.24 ;
     RECT  367.78 929.82 379.78 930.02 ;
     RECT  363 0 381 178 ;
     RECT  363 1622 381 1800 ;
     RECT  374.98 1308.66 381.22 1312.22 ;
     RECT  372.86 1331.34 381.5 1341.2 ;
     RECT  371.9 956.7 381.98 956.9 ;
     RECT  378.62 1356.96 383.14 1363.04 ;
     RECT  379.1 942.42 383.42 943.04 ;
     RECT  381.98 953.76 383.42 956.9 ;
     RECT  374.98 1289.76 383.9 1299.2 ;
     RECT  372.58 969.3 384.38 969.5 ;
     RECT  373.54 978.54 384.38 978.74 ;
     RECT  379.19 219.14 384.81 884.24 ;
     RECT  384.38 969.3 384.86 978.74 ;
     RECT  383.42 942.42 385.34 956.9 ;
     RECT  384.86 968.46 385.34 978.74 ;
     RECT  244.22 1449.32 385.34 1468.84 ;
     RECT  376.42 1126.8 385.82 1255.52 ;
     RECT  383.9 1289.76 385.82 1299.62 ;
     RECT  381.22 1308.66 385.82 1310.54 ;
     RECT  383.14 1359.06 386.3 1363.04 ;
     RECT  376.7 1371.66 386.3 1389.08 ;
     RECT  386.3 1359.06 386.78 1389.08 ;
     RECT  385.34 942.42 386.98 978.74 ;
     RECT  385.82 1289.76 387.74 1310.54 ;
     RECT  384.81 381.26 387.94 575.5 ;
     RECT  376.42 1006.26 388.22 1114.4 ;
     RECT  385.34 1449.32 388.22 1475.18 ;
     RECT  388.22 1006.26 388.7 1116.92 ;
     RECT  385.82 1126.8 388.7 1256.36 ;
     RECT  381.98 930.66 388.9 930.86 ;
     RECT  374.3 1272.96 389.18 1275.68 ;
     RECT  387.74 1288.92 389.18 1310.54 ;
     RECT  382.94 1319.58 389.38 1319.78 ;
     RECT  388.22 1445.16 389.38 1475.18 ;
     RECT  389.38 1445.16 389.66 1468.84 ;
     RECT  372.1 991.98 390.14 994.7 ;
     RECT  388.7 1006.26 390.14 1256.36 ;
     RECT  390.14 991.98 390.34 1256.36 ;
     RECT  381.5 1331.34 390.34 1346.66 ;
     RECT  389.18 1272.96 390.62 1310.54 ;
     RECT  390.34 1333.86 390.62 1346.66 ;
     RECT  390.34 1103.28 391.1 1256.36 ;
     RECT  391.1 1103.28 391.3 1260.56 ;
     RECT  390.62 1333.86 392.06 1350.02 ;
     RECT  386.78 1359.06 392.06 1389.5 ;
     RECT  392.06 1333.86 392.26 1389.5 ;
     RECT  392.26 1375.86 393.5 1389.5 ;
     RECT  392.26 1333.86 393.7 1364.72 ;
     RECT  393.7 1349.82 394.66 1364.72 ;
     RECT  393.7 1333.86 396.1 1335.32 ;
     RECT  391.3 1208.7 397.34 1260.56 ;
     RECT  390.62 1272.96 397.34 1316 ;
     RECT  397.34 1208.7 397.54 1316 ;
     RECT  397.54 1240.62 397.82 1316 ;
     RECT  389.66 1438.44 397.82 1468.84 ;
     RECT  386.98 942.42 398.3 956.9 ;
     RECT  390.34 991.98 398.78 1092.98 ;
     RECT  391.3 1103.28 398.78 1200.08 ;
     RECT  398.3 942.42 399.26 957.32 ;
     RECT  386.98 968.46 399.26 978.74 ;
     RECT  384.86 1406.1 399.26 1406.3 ;
     RECT  398.78 991.98 399.74 1200.08 ;
     RECT  397.54 1208.7 399.74 1229.06 ;
     RECT  399.26 942.42 400.22 978.74 ;
     RECT  400.22 938.64 401.66 978.74 ;
     RECT  399.74 991.98 401.86 1229.06 ;
     RECT  397.82 1436.76 402.34 1468.84 ;
     RECT  393.5 1375.86 402.82 1392.44 ;
     RECT  394.66 1359.06 403.1 1364.72 ;
     RECT  399.26 1406.1 403.3 1410.5 ;
     RECT  387.94 404.78 403.58 575.5 ;
     RECT  397.82 1240.62 403.78 1318.94 ;
     RECT  403.58 404.78 404.06 576.76 ;
     RECT  401.66 933.6 404.06 978.74 ;
     RECT  402.82 1375.86 404.26 1392.02 ;
     RECT  403.3 1407.36 406.46 1410.5 ;
     RECT  405.5 1422.48 406.46 1422.68 ;
     RECT  404.06 933.6 406.66 979.58 ;
     RECT  402.34 1438.44 406.66 1468.84 ;
     RECT  406.46 1407.36 407.9 1413.86 ;
     RECT  406.46 1422.48 407.9 1427.3 ;
     RECT  407.9 1407.36 408.1 1427.3 ;
     RECT  401.86 991.98 408.58 1227.8 ;
     RECT  396.1 1333.86 408.58 1334.06 ;
     RECT  406.66 933.6 409.06 978.74 ;
     RECT  384.81 852.92 410.3 884.24 ;
     RECT  409.06 934.44 410.5 978.74 ;
     RECT  403.1 1359.06 411.74 1365.14 ;
     RECT  410.5 939.06 411.94 968.66 ;
     RECT  411.94 950.4 412.42 968.66 ;
     RECT  403.78 1240.62 412.9 1309.28 ;
     RECT  410.5 978.54 413.38 978.74 ;
     RECT  403.78 1318.74 413.66 1318.94 ;
     RECT  411.74 1359.06 413.66 1365.56 ;
     RECT  404.26 1377.96 413.66 1392.02 ;
     RECT  413.66 1359.06 414.14 1392.02 ;
     RECT  408.1 1407.36 414.14 1414.7 ;
     RECT  381 1622 414.14 1870 ;
     RECT  412.42 968.46 414.34 968.66 ;
     RECT  394.66 1349.82 415.58 1350.02 ;
     RECT  414.14 1359.06 415.58 1414.7 ;
     RECT  408.1 1427.1 415.58 1427.3 ;
     RECT  406.66 1438.44 415.58 1438.64 ;
     RECT  415.58 1427.1 416.54 1438.64 ;
     RECT  415.58 1349.82 416.74 1414.7 ;
     RECT  408.58 991.98 417.22 1198.82 ;
     RECT  412.9 1263.72 417.22 1309.28 ;
     RECT  416.74 1377.96 417.22 1414.7 ;
     RECT  414.14 1620.68 417.5 1870 ;
     RECT  417.22 1409.04 417.7 1414.7 ;
     RECT  408.58 1208.7 419.14 1227.8 ;
     RECT  417.22 1263.72 419.14 1263.92 ;
     RECT  417.7 1409.88 419.42 1414.7 ;
     RECT  416.54 1425.84 419.42 1438.64 ;
     RECT  411.94 939.06 420.58 939.26 ;
     RECT  417.22 1003.74 420.58 1198.82 ;
     RECT  413.66 1318.74 420.86 1327.34 ;
     RECT  412.42 950.4 421.34 956.9 ;
     RECT  419.14 1225.5 421.34 1227.8 ;
     RECT  412.9 1240.62 421.34 1253.84 ;
     RECT  416.74 1349.82 421.34 1366.4 ;
     RECT  404.06 404.36 421.82 576.76 ;
     RECT  421.34 949.56 421.82 956.9 ;
     RECT  421.34 1225.5 421.82 1253.84 ;
     RECT  417.5 926.46 422.5 926.66 ;
     RECT  420.58 1006.68 422.78 1198.82 ;
     RECT  419.14 1208.7 422.78 1215.2 ;
     RECT  419.42 1409.88 423.74 1438.64 ;
     RECT  423.74 968.46 424.22 968.66 ;
     RECT  424.22 968.46 424.7 976.22 ;
     RECT  421.34 1346.46 424.7 1366.4 ;
     RECT  417.22 1272.96 425.18 1309.28 ;
     RECT  420.86 1318.74 425.18 1329.44 ;
     RECT  424.7 1338.9 425.18 1366.4 ;
     RECT  421.82 949.14 425.66 956.9 ;
     RECT  424.7 968.04 425.66 976.64 ;
     RECT  417.22 991.98 427.1 994.7 ;
     RECT  417.22 1377.96 427.3 1400.42 ;
     RECT  425.18 1272.96 427.58 1366.4 ;
     RECT  427.3 1377.96 427.58 1381.52 ;
     RECT  423.74 1409.88 427.58 1440.74 ;
     RECT  406.66 1449.32 427.58 1468.84 ;
     RECT  421.82 1225.5 428.06 1263.5 ;
     RECT  422.78 1006.68 428.54 1215.2 ;
     RECT  428.06 1225.5 428.54 1263.92 ;
     RECT  427.58 1272.96 428.54 1381.52 ;
     RECT  425.66 949.14 429.02 976.64 ;
     RECT  427.1 989.04 429.02 994.7 ;
     RECT  428.54 1006.68 429.02 1381.52 ;
     RECT  429.02 949.14 429.5 994.7 ;
     RECT  429.02 1006.26 429.5 1381.52 ;
     RECT  427.3 1390.98 430.18 1400.42 ;
     RECT  429.02 926.04 430.46 926.24 ;
     RECT  429.5 949.14 430.94 1381.52 ;
     RECT  430.46 921.42 432.86 926.24 ;
     RECT  432.86 914.7 433.82 926.24 ;
     RECT  430.94 942.84 434.98 1381.52 ;
     RECT  434.98 942.84 436.7 1225.7 ;
     RECT  430.18 1391.4 436.7 1400.42 ;
     RECT  427.58 1409.88 436.7 1468.84 ;
     RECT  434.98 1237.26 437.18 1381.52 ;
     RECT  387.94 381.26 437.66 395.32 ;
     RECT  421.82 404.36 437.66 577.18 ;
     RECT  436.7 940.74 437.66 1225.7 ;
     RECT  437.18 1237.26 438.34 1382.36 ;
     RECT  436.7 1391.4 438.34 1468.84 ;
     RECT  438.34 1343.94 439.78 1382.36 ;
     RECT  438.34 1237.26 440.26 1335.32 ;
     RECT  437.66 938.64 440.54 1225.7 ;
     RECT  433.82 914.7 441.02 926.66 ;
     RECT  440.54 938.22 441.02 1225.7 ;
     RECT  441.02 914.7 442.66 1225.7 ;
     RECT  438.34 1391.82 442.66 1468.84 ;
     RECT  442.66 914.7 443.62 995.96 ;
     RECT  439.78 1346.46 443.62 1382.36 ;
     RECT  442.66 1392.24 444.58 1468.84 ;
     RECT  443.62 1346.46 446.02 1380.68 ;
     RECT  442.66 1006.26 446.5 1225.7 ;
     RECT  444.58 1417.44 446.5 1468.84 ;
     RECT  444.58 1392.24 448.42 1407.56 ;
     RECT  446.02 1354.44 448.9 1380.68 ;
     RECT  446.5 1018.44 449.38 1225.7 ;
     RECT  448.9 1354.44 450.34 1377.74 ;
     RECT  440.26 1237.26 450.62 1311.8 ;
     RECT  440.26 1323.78 450.62 1335.32 ;
     RECT  449.38 1018.44 450.82 1215.2 ;
     RECT  450.62 1237.26 450.82 1335.32 ;
     RECT  381 -70 451 178 ;
     RECT  417.5 1620.26 451 1870 ;
     RECT  443.62 978.54 451.1 995.96 ;
     RECT  450.82 1320 451.78 1335.32 ;
     RECT  443.62 914.7 452.06 969.08 ;
     RECT  451.1 978.54 452.06 996.38 ;
     RECT  450.34 1354.44 452.26 1373.12 ;
     RECT  448.42 1398.96 452.26 1407.56 ;
     RECT  450.82 1028.1 452.74 1215.2 ;
     RECT  451.78 1320 452.74 1329.86 ;
     RECT  446.5 1417.86 453.22 1468.84 ;
     RECT  452.26 1399.38 453.7 1407.56 ;
     RECT  446.5 1006.26 455.9 1006.46 ;
     RECT  450.82 1018.44 455.9 1019.06 ;
     RECT  452.26 1354.44 456.1 1365.14 ;
     RECT  453.7 1403.58 457.34 1407.56 ;
     RECT  453.22 1417.86 457.34 1422.26 ;
     RECT  455.9 1006.26 457.54 1019.06 ;
     RECT  450.82 1237.26 457.54 1309.28 ;
     RECT  457.54 1237.26 458.02 1263.92 ;
     RECT  452.06 914.7 459.26 996.38 ;
     RECT  457.54 1006.26 459.26 1006.46 ;
     RECT  457.34 1403.58 460.42 1422.26 ;
     RECT  452.74 1207.02 460.7 1215.2 ;
     RECT  449.38 1225.08 460.7 1225.7 ;
     RECT  457.54 1018.44 461.18 1019.06 ;
     RECT  452.74 1028.1 461.18 1195.04 ;
     RECT  459.26 914.7 461.38 1006.46 ;
     RECT  460.7 1207.02 461.38 1225.7 ;
     RECT  410.3 852.92 461.66 889.7 ;
     RECT  381.5 905.46 461.66 905.66 ;
     RECT  457.54 1272.96 461.86 1309.28 ;
     RECT  461.66 852.92 462.14 905.66 ;
     RECT  461.38 914.7 462.14 994.7 ;
     RECT  461.38 1207.02 462.14 1215.2 ;
     RECT  462.14 852.92 463.3 994.7 ;
     RECT  460.42 1403.58 463.3 1418.06 ;
     RECT  463.3 1403.58 464.54 1415.12 ;
     RECT  463.3 915.54 464.74 994.7 ;
     RECT  461.86 1272.96 464.74 1293.74 ;
     RECT  461.18 1018.44 465.22 1195.04 ;
     RECT  461.38 1224.66 465.22 1225.7 ;
     RECT  461.86 1308.66 465.98 1309.28 ;
     RECT  452.74 1320 465.98 1326.92 ;
     RECT  464.54 1395.18 465.98 1415.12 ;
     RECT  456.1 1354.44 466.66 1354.64 ;
     RECT  458.02 1237.26 466.94 1262.66 ;
     RECT  464.74 915.54 467.14 939.26 ;
     RECT  464.74 948.3 467.14 994.7 ;
     RECT  464.74 1272.96 467.14 1289.96 ;
     RECT  466.94 1236 467.62 1262.66 ;
     RECT  465.98 1308.66 468.1 1326.92 ;
     RECT  467.14 915.54 468.58 936.74 ;
     RECT  451 0 469 178 ;
     RECT  451 1620.26 469 1800 ;
     RECT  467.14 1286.4 469.06 1289.96 ;
     RECT  467.62 1236 469.54 1260.14 ;
     RECT  465.22 1018.44 470.5 1193.78 ;
     RECT  469.06 1286.4 470.5 1287.44 ;
     RECT  467.42 1349.82 470.5 1350.02 ;
     RECT  465.98 1387.2 470.5 1415.12 ;
     RECT  467.14 948.3 470.98 961.1 ;
     RECT  468.1 1308.66 470.98 1319.36 ;
     RECT  462.14 1206.6 471.46 1215.2 ;
     RECT  465.22 1224.66 471.46 1225.28 ;
     RECT  453.22 1431.3 471.46 1468.84 ;
     RECT  469.54 1236 471.94 1258.46 ;
     RECT  470.5 1387.2 471.94 1387.4 ;
     RECT  470.5 1403.58 471.94 1415.12 ;
     RECT  471.94 1410.3 472.9 1410.5 ;
     RECT  471.46 1209.96 473.18 1215.2 ;
     RECT  471.94 1243.98 473.38 1258.46 ;
     RECT  467.14 970.14 474.14 994.7 ;
     RECT  461.38 1006.26 474.14 1006.46 ;
     RECT  474.14 970.14 474.62 1006.46 ;
     RECT  473.18 1209.96 474.82 1223.6 ;
     RECT  471.46 1431.3 475.3 1449.94 ;
     RECT  475.3 1431.3 475.78 1440.74 ;
     RECT  475.78 1440.54 476.26 1440.74 ;
     RECT  468.58 918.06 476.54 936.74 ;
     RECT  470.98 949.14 476.54 961.1 ;
     RECT  470.5 1028.1 476.54 1193.78 ;
     RECT  470.98 1319.16 476.74 1319.36 ;
     RECT  476.54 949.14 477.5 961.52 ;
     RECT  474.62 970.14 477.5 1016.96 ;
     RECT  476.54 918.06 477.7 940.1 ;
     RECT  437.66 381.26 477.98 577.18 ;
     RECT  477.5 949.14 479.9 1016.96 ;
     RECT  476.54 1028.1 479.9 1196.72 ;
     RECT  470.98 1308.66 480.1 1309.28 ;
     RECT  463.3 852.92 481.82 905.66 ;
     RECT  477.7 918.48 481.82 940.1 ;
     RECT  479.9 949.14 481.82 1196.72 ;
     RECT  481.82 918.48 482.5 1196.72 ;
     RECT  394.46 348.92 482.78 349.12 ;
     RECT  482.5 918.9 483.74 1196.72 ;
     RECT  473.38 1243.98 483.74 1257.62 ;
     RECT  483.74 1236.42 484.9 1257.62 ;
     RECT  480.1 1309.08 484.9 1309.28 ;
     RECT  467.14 1272.96 485.86 1274.42 ;
     RECT  484.9 1243.98 489.7 1257.62 ;
     RECT  475.78 1431.3 490.18 1431.5 ;
     RECT  489.7 1243.98 490.66 1244.18 ;
     RECT  485.86 1274.22 491.14 1274.42 ;
     RECT  489.7 1257.42 491.62 1257.62 ;
     RECT  483.74 918.9 492.38 1197.14 ;
     RECT  474.82 1209.96 492.38 1219.82 ;
     RECT  470.5 1286.4 492.38 1286.6 ;
     RECT  492.38 918.9 492.86 1197.6 ;
     RECT  492.38 1280.56 495.94 1286.6 ;
     RECT  495.74 1238.98 496.22 1239.18 ;
     RECT  497.66 1404.88 498.14 1405.08 ;
     RECT  496.22 1236.46 499.58 1239.18 ;
     RECT  499.58 1265.02 500.06 1265.22 ;
     RECT  477.98 381.26 500.54 577.6 ;
     RECT  384.81 587.06 500.54 592.3 ;
     RECT  499.1 1352.38 500.54 1352.58 ;
     RECT  475.3 1449.32 501.5 1449.94 ;
     RECT  499.58 1236.46 502.46 1244.64 ;
     RECT  501.5 1306.18 502.46 1306.38 ;
     RECT  490.46 1424.62 502.46 1424.82 ;
     RECT  496.7 1435.96 502.46 1436.16 ;
     RECT  500.54 1349.86 503.62 1352.58 ;
     RECT  500.06 1265.02 503.9 1267.32 ;
     RECT  501.98 1296.1 504.38 1296.3 ;
     RECT  502.46 1236.46 504.58 1250.94 ;
     RECT  502.46 1424.62 504.58 1436.16 ;
     RECT  502.46 1306.18 504.86 1309.74 ;
     RECT  492.86 915.12 505.34 1197.6 ;
     RECT  495.94 1280.56 505.82 1280.76 ;
     RECT  504.38 1291.9 505.82 1296.3 ;
     RECT  490.46 1375.06 506.02 1375.26 ;
     RECT  503.9 1265.02 506.3 1269.42 ;
     RECT  505.82 1280.56 506.3 1296.3 ;
     RECT  505.34 915.12 507.26 1198.44 ;
     RECT  492.38 1209.96 507.26 1224.48 ;
     RECT  504.58 1236.46 507.26 1243.38 ;
     RECT  506.3 1263.76 507.26 1296.3 ;
     RECT  504.86 1306.18 508.22 1311.42 ;
     RECT  504.58 1435.54 508.22 1436.16 ;
     RECT  501.5 1446.88 508.22 1449.94 ;
     RECT  471.46 1459.4 508.22 1468.84 ;
     RECT  508.22 1306.18 509.18 1311.84 ;
     RECT  507.26 1260.82 509.38 1296.3 ;
     RECT  509.18 1306.18 509.38 1312.26 ;
     RECT  504.58 1424.62 509.38 1424.82 ;
     RECT  507.26 915.12 509.86 1243.38 ;
     RECT  507.74 1356.16 509.86 1356.36 ;
     RECT  507.74 1366.66 510.14 1366.86 ;
     RECT  509.38 1260.82 510.34 1292.1 ;
     RECT  510.34 1260.82 510.62 1274.88 ;
     RECT  510.34 1284.34 510.82 1292.1 ;
     RECT  510.82 1284.34 512.26 1284.54 ;
     RECT  509.86 919.32 513.02 1243.38 ;
     RECT  510.62 1258.3 513.02 1274.88 ;
     RECT  513.02 919.32 513.22 1274.88 ;
     RECT  498.14 1404.04 514.66 1405.08 ;
     RECT  510.62 1416.64 514.66 1418.1 ;
     RECT  405.02 327.5 515.19 327.7 ;
     RECT  482.78 341.78 515.19 349.12 ;
     RECT  500.54 381.26 515.19 592.3 ;
     RECT  384.81 601.34 515.19 842.62 ;
     RECT  481.82 852.08 515.19 905.66 ;
     RECT  316.81 1573.22 515.19 1583.08 ;
     RECT  510.14 1360.36 517.06 1366.86 ;
     RECT  509.38 1306.18 517.82 1311.84 ;
     RECT  508.22 1435.54 518.98 1449.94 ;
     RECT  513.22 1209.96 519.26 1274.88 ;
     RECT  519.26 1292.32 520.42 1292.52 ;
     RECT  517.82 1303.24 520.42 1311.84 ;
     RECT  515.19 215.36 520.7 905.66 ;
     RECT  513.22 919.32 520.7 1201.38 ;
     RECT  520.42 1309.54 520.7 1311.84 ;
     RECT  520.7 215.36 520.81 1201.38 ;
     RECT  515.19 1573.22 520.81 1583.92 ;
     RECT  508.22 1459.4 520.9 1469.76 ;
     RECT  519.26 1375.06 521.66 1375.26 ;
     RECT  520.7 1309.54 522.34 1312.26 ;
     RECT  495.74 1333.9 523.3 1334.1 ;
     RECT  514.66 1416.64 524.06 1417.68 ;
     RECT  518.98 1446.88 524.26 1449.94 ;
     RECT  515.9 1346.08 525.22 1346.28 ;
     RECT  521.66 1375.06 525.7 1381.14 ;
     RECT  519.26 1209.96 526.18 1281.18 ;
     RECT  524.06 1416.64 526.46 1424.82 ;
     RECT  526.18 1209.96 526.66 1244.22 ;
     RECT  517.82 1401.52 528.58 1401.72 ;
     RECT  526.66 1209.96 529.06 1242.96 ;
     RECT  526.18 1258.3 529.06 1281.18 ;
     RECT  520.81 601.34 529.54 1201.38 ;
     RECT  525.7 1375.9 530.78 1381.14 ;
     RECT  529.54 1201.18 530.98 1201.38 ;
     RECT  529.06 1209.96 530.98 1241.7 ;
     RECT  517.06 1360.36 530.98 1360.56 ;
     RECT  526.46 1413.7 531.94 1424.82 ;
     RECT  529.06 1258.3 532.42 1280.76 ;
     RECT  530.98 1209.96 533.38 1219.82 ;
     RECT  532.42 1258.3 533.38 1274.88 ;
     RECT  533.38 1212.48 533.86 1219.82 ;
     RECT  531.94 1413.7 534.34 1422.3 ;
     RECT  533.86 1212.48 534.82 1215.2 ;
     RECT  529.54 601.34 535.78 1192.52 ;
     RECT  533.38 1258.3 535.78 1274.46 ;
     RECT  534.82 1212.48 536.26 1214.78 ;
     RECT  535.78 1258.3 536.74 1272.36 ;
     RECT  530.78 1375.9 536.74 1383.24 ;
     RECT  534.34 1413.7 537.5 1413.9 ;
     RECT  530.98 1230.16 537.7 1241.7 ;
     RECT  536.74 1258.3 537.7 1269.84 ;
     RECT  536.74 1383.04 537.7 1383.24 ;
     RECT  522.34 1309.54 538.46 1309.74 ;
     RECT  520.9 1459.4 538.46 1468.84 ;
     RECT  469 -70 539 178 ;
     RECT  469 1620.26 539 1870 ;
     RECT  538.46 1309.54 541.34 1318.14 ;
     RECT  537.5 1291.06 541.82 1291.26 ;
     RECT  539.9 1341.46 541.82 1341.66 ;
     RECT  541.34 1201.18 542.3 1201.38 ;
     RECT  541.34 1309.54 542.3 1318.56 ;
     RECT  524.26 1449.32 542.3 1449.94 ;
     RECT  537.5 1409.92 542.78 1413.9 ;
     RECT  541.82 1341.46 543.26 1345.02 ;
     RECT  542.78 1401.94 543.46 1421.04 ;
     RECT  542.3 1197.4 545.38 1201.38 ;
     RECT  541.82 1287.28 546.62 1291.26 ;
     RECT  542.3 1304.08 546.62 1318.98 ;
     RECT  539.9 1364.14 546.62 1364.34 ;
     RECT  546.62 1287.28 546.82 1318.98 ;
     RECT  520.81 1573.22 546.82 1583.08 ;
     RECT  536.26 1212.48 547.3 1212.68 ;
     RECT  538.46 1459.4 548.26 1477.32 ;
     RECT  546.82 1287.28 548.74 1318.56 ;
     RECT  537.7 1265.86 549.02 1269.84 ;
     RECT  543.26 1341.46 549.02 1352.58 ;
     RECT  549.02 1265.44 549.22 1269.84 ;
     RECT  520.81 381.26 549.98 592.3 ;
     RECT  549.02 1337.68 549.98 1352.58 ;
     RECT  549.98 1337.26 550.46 1352.58 ;
     RECT  546.62 1364.14 550.46 1364.76 ;
     RECT  550.46 1337.26 551.9 1364.76 ;
     RECT  548.74 1287.28 552.1 1318.14 ;
     RECT  543.46 1401.94 552.38 1405.92 ;
     RECT  542.3 1443.52 553.54 1449.94 ;
     RECT  543.46 1417.06 553.82 1421.04 ;
     RECT  537.7 1230.16 554.3 1239.18 ;
     RECT  553.82 1417.06 554.3 1427.76 ;
     RECT  551.9 1331.38 555.46 1364.76 ;
     RECT  554.3 1417.06 555.74 1428.6 ;
     RECT  552.38 1393.96 556.42 1405.92 ;
     RECT  539 0 557 178 ;
     RECT  539 1620.26 557 1800 ;
     RECT  545.38 1197.4 557.18 1197.6 ;
     RECT  551.9 1208.74 557.18 1208.94 ;
     RECT  549.22 1269.22 557.18 1269.84 ;
     RECT  552.1 1287.28 558.34 1314.78 ;
     RECT  557.18 1208.74 558.82 1216.08 ;
     RECT  553.82 1254.52 559.1 1254.72 ;
     RECT  557.18 1269.22 559.1 1273.62 ;
     RECT  557.18 1196.98 559.3 1197.6 ;
     RECT  556.42 1393.96 559.78 1402.14 ;
     RECT  559.78 1401.94 561.22 1402.14 ;
     RECT  554.3 1230.16 562.94 1243.38 ;
     RECT  555.74 1417.06 563.14 1439.94 ;
     RECT  558.34 1290.64 563.62 1314.78 ;
     RECT  555.46 1344.82 564.38 1364.76 ;
     RECT  558.82 1208.74 564.58 1208.94 ;
     RECT  563.14 1417.06 566.3 1435.74 ;
     RECT  566.3 1412.86 566.5 1435.74 ;
     RECT  535.78 601.34 566.78 1186.22 ;
     RECT  564.38 1341.88 566.78 1364.76 ;
     RECT  564.38 1373.38 566.78 1373.58 ;
     RECT  559.58 1383.04 566.98 1383.24 ;
     RECT  563.62 1290.64 567.74 1295.46 ;
     RECT  563.62 1307.44 568.22 1314.78 ;
     RECT  568.22 1307.44 568.7 1316.04 ;
     RECT  559.1 1254.52 568.9 1273.62 ;
     RECT  566.78 601.34 569.18 1186.26 ;
     RECT  559.3 1197.4 569.18 1197.6 ;
     RECT  568.7 1307.44 569.66 1316.46 ;
     RECT  568.9 1261.24 570.14 1273.62 ;
     RECT  569.18 601.34 570.34 1197.6 ;
     RECT  569.66 1307.44 570.82 1323.6 ;
     RECT  562.94 1223.86 571.78 1243.38 ;
     RECT  570.14 1261.24 571.78 1274.46 ;
     RECT  566.5 1412.86 571.78 1432.38 ;
     RECT  570.34 601.34 572.74 1192.14 ;
     RECT  567.74 1286.44 572.74 1295.46 ;
     RECT  566.78 1341.88 572.74 1373.58 ;
     RECT  571.78 1223.86 573.02 1236.24 ;
     RECT  573.02 1217.14 573.22 1236.24 ;
     RECT  572.74 1289.38 575.14 1295.46 ;
     RECT  572.74 1341.88 575.9 1352.58 ;
     RECT  572.74 1163.76 576.1 1192.14 ;
     RECT  571.78 1262.08 577.54 1273.62 ;
     RECT  575.9 1341.46 577.82 1352.58 ;
     RECT  577.54 1269.22 578.5 1273.62 ;
     RECT  576.1 1186.9 578.98 1192.14 ;
     RECT  570.82 1307.44 579.46 1318.98 ;
     RECT  577.82 1338.52 580.9 1352.58 ;
     RECT  578.98 1186.9 581.38 1187.1 ;
     RECT  573.22 1217.14 581.86 1235.4 ;
     RECT  576.38 1298.2 582.34 1298.4 ;
     RECT  576.38 1327.6 582.34 1327.8 ;
     RECT  576.1 1163.76 582.82 1177.82 ;
     RECT  581.86 1217.14 582.82 1217.34 ;
     RECT  575.14 1289.38 583.1 1289.58 ;
     RECT  520.81 255.26 583.19 255.46 ;
     RECT  570.62 269.96 583.19 270.16 ;
     RECT  520.81 327.5 583.19 327.7 ;
     RECT  520.81 341.78 583.19 349.12 ;
     RECT  549.98 380.84 583.19 592.3 ;
     RECT  572.74 601.34 583.19 1154.72 ;
     RECT  546.82 1573.22 583.19 1579.3 ;
     RECT  571.78 1417.06 583.3 1432.38 ;
     RECT  583.1 1283.92 584.26 1289.58 ;
     RECT  579.46 1307.44 584.74 1314.36 ;
     RECT  572.74 1364.56 584.74 1373.58 ;
     RECT  584.74 1307.44 585.98 1307.64 ;
     RECT  582.62 1256.62 586.66 1256.82 ;
     RECT  578.5 1269.22 586.94 1270.26 ;
     RECT  585.5 1330.12 587.14 1330.32 ;
     RECT  585.98 1306.18 587.62 1307.64 ;
     RECT  580.9 1339.36 587.62 1352.58 ;
     RECT  586.94 1259.98 587.9 1260.18 ;
     RECT  586.94 1269.22 587.9 1271.1 ;
     RECT  584.74 1373.38 587.9 1373.58 ;
     RECT  581.86 1226.8 588.1 1235.4 ;
     RECT  584.26 1289.38 588.1 1289.58 ;
     RECT  587.62 1307.44 588.1 1307.64 ;
     RECT  587.62 1339.36 588.1 1351.32 ;
     RECT  587.9 1373.38 588.1 1380.72 ;
     RECT  553.54 1449.32 588.38 1449.94 ;
     RECT  548.26 1459.4 588.38 1468.84 ;
     RECT  587.9 1259.98 588.58 1271.1 ;
     RECT  583.19 219.14 588.81 1154.72 ;
     RECT  583.19 1573.22 588.81 1580.14 ;
     RECT  584.74 1364.56 589.06 1364.76 ;
     RECT  582.82 1164.18 589.34 1177.82 ;
     RECT  588.86 1192.78 590.3 1192.98 ;
     RECT  588.1 1226.8 590.3 1229.52 ;
     RECT  589.34 1410.34 590.78 1410.54 ;
     RECT  588.38 1238.98 591.46 1241.7 ;
     RECT  590.3 1220.5 591.94 1229.52 ;
     RECT  588.81 601.34 592.42 1154.72 ;
     RECT  589.34 1164.18 592.7 1178.28 ;
     RECT  592.42 926.04 592.9 1150.52 ;
     RECT  587.9 1209.58 592.9 1209.78 ;
     RECT  588.58 1262.08 593.18 1271.1 ;
     RECT  583.3 1424.62 593.18 1432.38 ;
     RECT  592.9 927.3 593.38 1150.52 ;
     RECT  587.9 1320.46 593.66 1320.66 ;
     RECT  590.78 1409.5 593.66 1410.54 ;
     RECT  593.66 1409.5 593.86 1413.06 ;
     RECT  593.18 1422.1 594.14 1432.38 ;
     RECT  592.22 1293.58 594.62 1293.78 ;
     RECT  591.94 1220.5 595.1 1229.1 ;
     RECT  591.46 1238.98 595.3 1239.18 ;
     RECT  593.86 1409.92 595.3 1413.06 ;
     RECT  592.7 1390.18 595.58 1390.38 ;
     RECT  594.14 1421.68 596.06 1432.38 ;
     RECT  593.18 1262.08 597.02 1273.2 ;
     RECT  593.66 1311.64 597.02 1320.66 ;
     RECT  595.58 1390.18 597.5 1394.16 ;
     RECT  595.1 1216.72 598.18 1229.1 ;
     RECT  597.02 1258.72 598.46 1273.2 ;
     RECT  594.62 1293.58 599.42 1295.04 ;
     RECT  588.1 1339.36 599.42 1339.56 ;
     RECT  588.1 1351.12 599.42 1351.32 ;
     RECT  592.7 1164.18 599.9 1179.12 ;
     RECT  590.3 1187.74 599.9 1192.98 ;
     RECT  597.02 1309.12 600.58 1320.66 ;
     RECT  599.42 1292.74 600.86 1295.04 ;
     RECT  599.42 1337.68 601.54 1339.56 ;
     RECT  597.5 1390.18 601.54 1397.94 ;
     RECT  601.54 1337.68 602.02 1337.88 ;
     RECT  592.42 601.34 602.78 916.16 ;
     RECT  593.38 927.3 602.78 1145.06 ;
     RECT  598.46 1251.58 602.98 1273.2 ;
     RECT  596.06 1421.68 603.74 1439.94 ;
     RECT  588.38 1449.32 603.74 1468.84 ;
     RECT  602.78 601.34 604.7 1145.06 ;
     RECT  603.74 1421.68 604.9 1468.84 ;
     RECT  600.86 1291.9 605.18 1295.04 ;
     RECT  595.3 1412.02 605.66 1413.06 ;
     RECT  604.9 1421.68 605.66 1449.94 ;
     RECT  599.9 1164.18 606.14 1192.98 ;
     RECT  604.9 1459.4 606.14 1468.84 ;
     RECT  598.18 1216.72 607.3 1224.48 ;
     RECT  606.14 1164.18 607.58 1198.86 ;
     RECT  588.1 1373.8 608.54 1380.72 ;
     RECT  601.54 1390.18 608.54 1390.38 ;
     RECT  599.42 1351.12 609.02 1356.36 ;
     RECT  605.66 1412.02 609.02 1449.94 ;
     RECT  605.18 1280.14 609.98 1281.18 ;
     RECT  605.18 1291.06 609.98 1295.04 ;
     RECT  602.98 1251.58 611.42 1269.84 ;
     RECT  609.02 1348.6 611.42 1356.36 ;
     RECT  608.54 1373.8 611.42 1390.38 ;
     RECT  609.02 1406.14 611.62 1449.94 ;
     RECT  588.81 341.78 611.9 349.12 ;
     RECT  611.42 1251.58 612.38 1271.52 ;
     RECT  609.98 1280.14 612.38 1295.04 ;
     RECT  607.58 1164.18 612.58 1201.8 ;
     RECT  612.38 1251.58 613.06 1295.04 ;
     RECT  611.42 1348.6 613.82 1356.78 ;
     RECT  611.42 1373.8 614.78 1396.68 ;
     RECT  611.62 1410.34 614.98 1449.94 ;
     RECT  588.81 380.84 615.26 592.3 ;
     RECT  604.7 601.34 615.26 1151.82 ;
     RECT  612.58 1170.94 615.94 1201.8 ;
     RECT  614.78 1367.08 616.42 1396.68 ;
     RECT  600.58 1311.22 616.7 1320.66 ;
     RECT  616.7 1303.66 616.9 1320.66 ;
     RECT  613.82 1343.56 617.18 1356.78 ;
     RECT  606.14 1459.4 618.82 1477.32 ;
     RECT  615.26 380.84 619.1 1151.82 ;
     RECT  616.9 1304.08 619.3 1320.66 ;
     RECT  617.18 1337.68 620.06 1356.78 ;
     RECT  614.98 1420.42 620.26 1449.94 ;
     RECT  615.94 1170.94 620.74 1186.26 ;
     RECT  617.18 1238.14 620.74 1238.34 ;
     RECT  619.1 380.84 621.98 1156.02 ;
     RECT  620.06 1333.9 621.98 1356.78 ;
     RECT  621.98 1331.8 622.46 1356.78 ;
     RECT  620.74 1175.14 622.66 1186.26 ;
     RECT  621.98 380.84 622.94 1156.44 ;
     RECT  619.3 1311.22 623.14 1320.66 ;
     RECT  622.46 1330.54 623.14 1356.78 ;
     RECT  623.14 1330.54 623.62 1343.76 ;
     RECT  615.94 1197.82 624.38 1201.8 ;
     RECT  613.06 1251.58 624.38 1281.18 ;
     RECT  613.06 1291.48 624.38 1295.04 ;
     RECT  614.98 1410.34 625.06 1410.54 ;
     RECT  622.94 380.84 625.54 1160.22 ;
     RECT  624.38 1251.58 625.54 1295.04 ;
     RECT  616.42 1367.08 626.5 1382.82 ;
     RECT  625.54 1292.74 626.98 1295.04 ;
     RECT  557 -70 627 178 ;
     RECT  557 1620.26 627 1870 ;
     RECT  622.66 1175.14 627.46 1184.16 ;
     RECT  626.98 1293.58 627.94 1295.04 ;
     RECT  623.14 1356.58 627.94 1356.78 ;
     RECT  625.54 1251.58 628.42 1279.08 ;
     RECT  626.5 1367.08 628.42 1379.46 ;
     RECT  623.14 1311.22 628.7 1311.42 ;
     RECT  628.42 1367.08 628.7 1371.9 ;
     RECT  628.7 1306.18 629.38 1311.42 ;
     RECT  628.42 1251.58 629.86 1276.98 ;
     RECT  628.7 1360.78 629.86 1371.9 ;
     RECT  629.38 1306.18 630.34 1306.38 ;
     RECT  620.26 1420.42 630.82 1432.38 ;
     RECT  623.62 1331.38 631.3 1343.76 ;
     RECT  627.94 1293.58 632.26 1293.78 ;
     RECT  629.86 1371.7 632.74 1371.9 ;
     RECT  627.46 1175.14 633.7 1182.06 ;
     RECT  623.14 1320.46 633.7 1320.66 ;
     RECT  631.3 1331.38 633.7 1334.1 ;
     RECT  624.38 1197.4 633.98 1201.8 ;
     RECT  620.26 1447.72 634.66 1449.94 ;
     RECT  633.98 1195.72 635.14 1201.8 ;
     RECT  635.14 1195.72 635.62 1198.86 ;
     RECT  631.58 1405.72 635.62 1405.92 ;
     RECT  631.3 1343.56 635.9 1343.76 ;
     RECT  629.86 1253.68 636.1 1276.98 ;
     RECT  635.9 1343.56 636.1 1346.28 ;
     RECT  630.82 1422.1 636.1 1432.38 ;
     RECT  636.1 1276.78 636.58 1276.98 ;
     RECT  633.7 1333.9 637.06 1334.1 ;
     RECT  636.1 1422.1 637.06 1422.3 ;
     RECT  633.5 1231.42 637.82 1231.62 ;
     RECT  616.42 1396.48 637.82 1396.68 ;
     RECT  636.1 1431.76 637.82 1432.38 ;
     RECT  633.7 1175.14 638.02 1181.22 ;
     RECT  629.86 1360.78 638.02 1360.98 ;
     RECT  637.82 1230.16 638.3 1235.82 ;
     RECT  637.82 1396.48 638.3 1403.82 ;
     RECT  636.1 1346.08 638.5 1346.28 ;
     RECT  630.62 1211.68 638.78 1211.88 ;
     RECT  638.3 1229.74 638.78 1235.82 ;
     RECT  638.3 1393.96 639.46 1403.82 ;
     RECT  638.78 1211.68 639.74 1213.14 ;
     RECT  639.26 1290.64 639.74 1291.26 ;
     RECT  639.46 1396.06 639.94 1397.94 ;
     RECT  639.74 1211.68 640.22 1218.18 ;
     RECT  638.78 1229.32 640.22 1235.82 ;
     RECT  640.22 1211.68 640.7 1235.82 ;
     RECT  639.74 1290.22 641.66 1291.26 ;
     RECT  640.7 1211.68 641.86 1240.86 ;
     RECT  641.86 1211.68 642.14 1240.02 ;
     RECT  638.02 1181.02 642.62 1181.22 ;
     RECT  641.18 1281.4 642.62 1281.6 ;
     RECT  641.66 1290.22 642.62 1293.78 ;
     RECT  634.66 1449.32 643.1 1449.94 ;
     RECT  618.82 1459.4 643.1 1468.84 ;
     RECT  643.1 1311.64 643.58 1311.84 ;
     RECT  625.54 380.84 644.06 1156.44 ;
     RECT  641.18 1171.36 644.06 1171.56 ;
     RECT  642.62 1281.4 644.06 1293.78 ;
     RECT  642.62 1181.02 644.26 1183.74 ;
     RECT  627 0 645 178 ;
     RECT  627 1620.26 645 1800 ;
     RECT  642.14 1210.84 646.18 1240.02 ;
     RECT  644.06 1281.4 646.18 1299.66 ;
     RECT  642.14 1350.28 646.18 1350.48 ;
     RECT  643.1 1449.32 646.66 1468.84 ;
     RECT  636.1 1253.68 646.94 1268.16 ;
     RECT  637.82 1431.76 647.14 1436.16 ;
     RECT  635.62 1198.66 647.62 1198.86 ;
     RECT  643.58 1311.64 647.9 1318.98 ;
     RECT  640.22 1416.22 647.9 1416.42 ;
     RECT  646.94 1253.68 648.1 1269.84 ;
     RECT  647.9 1303.24 648.58 1318.98 ;
     RECT  644.06 380.84 648.86 1171.56 ;
     RECT  639.74 1367.5 648.86 1367.7 ;
     RECT  648.86 380.84 649.06 1179.12 ;
     RECT  648.86 1367.5 649.34 1371.48 ;
     RECT  647.9 1416.22 649.34 1417.26 ;
     RECT  648.1 1253.68 649.82 1268.16 ;
     RECT  649.34 1364.14 649.82 1371.48 ;
     RECT  646.18 1212.94 650.02 1240.02 ;
     RECT  649.82 1249.9 650.98 1268.16 ;
     RECT  647.14 1432.18 651.46 1436.16 ;
     RECT  646.18 1281.4 651.74 1294.62 ;
     RECT  650.02 1212.94 651.94 1239.6 ;
     RECT  650.98 1253.68 651.94 1268.16 ;
     RECT  651.46 1432.18 651.94 1435.32 ;
     RECT  639.94 1396.48 652.42 1397.94 ;
     RECT  649.34 1412.02 652.42 1417.26 ;
     RECT  648.58 1303.24 652.9 1311.84 ;
     RECT  649.82 1363.72 653.66 1371.48 ;
     RECT  651.74 1279.72 655.78 1294.62 ;
     RECT  651.94 1257.88 656.74 1268.16 ;
     RECT  638.3 1477.96 656.74 1478.16 ;
     RECT  655.78 1284.76 657.22 1294.62 ;
     RECT  588.81 327.5 658.46 327.7 ;
     RECT  611.9 341.78 658.46 356.26 ;
     RECT  657.98 1328.86 658.94 1329.06 ;
     RECT  646.66 1449.32 658.94 1449.94 ;
     RECT  646.66 1459.4 658.94 1468.84 ;
     RECT  651.94 1215.88 659.14 1239.6 ;
     RECT  653.66 1363.72 659.14 1372.74 ;
     RECT  652.9 1307.44 659.62 1311.84 ;
     RECT  659.14 1367.5 660.1 1372.74 ;
     RECT  660.38 1204.96 661.34 1205.16 ;
     RECT  651.94 1432.18 661.34 1432.38 ;
     RECT  652.42 1412.02 661.54 1416.42 ;
     RECT  649.06 380.84 662.02 1163.16 ;
     RECT  659.14 1216.3 662.3 1239.6 ;
     RECT  657.22 1290.64 662.3 1294.62 ;
     RECT  659.62 1307.44 662.3 1307.64 ;
     RECT  658.94 1325.08 662.3 1329.06 ;
     RECT  649.06 1178.92 662.98 1179.12 ;
     RECT  656.54 1352.8 663.26 1353 ;
     RECT  661.34 1204.96 663.46 1205.58 ;
     RECT  662.3 1325.08 666.14 1332 ;
     RECT  662.3 1290.64 666.82 1307.64 ;
     RECT  662.02 380.84 667.3 1156.44 ;
     RECT  666.82 1290.64 667.58 1294.62 ;
     RECT  666.14 1324.66 669.02 1332 ;
     RECT  663.26 1346.5 669.02 1353 ;
     RECT  662.3 1216.3 669.7 1240.02 ;
     RECT  656.74 1258.3 669.98 1266.06 ;
     RECT  669.98 1251.16 670.18 1266.06 ;
     RECT  652.42 1396.48 670.18 1396.68 ;
     RECT  669.7 1216.3 671.62 1232.88 ;
     RECT  670.18 1251.16 671.62 1264.38 ;
     RECT  661.34 1432.18 671.62 1439.94 ;
     RECT  671.62 1256.2 673.06 1264.38 ;
     RECT  671.62 1432.18 673.06 1432.38 ;
     RECT  667.58 1288.54 673.82 1294.62 ;
     RECT  671.62 1216.3 674.02 1229.94 ;
     RECT  673.06 1256.2 674.02 1263.96 ;
     RECT  674.02 1221.34 674.5 1229.94 ;
     RECT  662.78 1189.84 674.78 1190.04 ;
     RECT  673.82 1282.24 674.78 1294.62 ;
     RECT  669.02 1324.66 674.78 1353 ;
     RECT  674.5 1221.34 674.98 1228.68 ;
     RECT  674.78 1319.2 674.98 1353 ;
     RECT  674.98 1319.2 675.46 1333.26 ;
     RECT  675.46 1319.2 675.94 1332.84 ;
     RECT  674.98 1346.5 676.42 1353 ;
     RECT  645 1620.26 677.86 1870 ;
     RECT  667.3 380.84 679.1 981.26 ;
     RECT  667.3 991.14 679.1 1156.44 ;
     RECT  674.78 1280.56 680.26 1294.62 ;
     RECT  680.26 1282.66 680.74 1294.62 ;
     RECT  676.42 1352.8 681.22 1353 ;
     RECT  658.94 1449.32 681.22 1468.84 ;
     RECT  674.02 1258.72 682.94 1263.96 ;
     RECT  679.1 380.84 683.14 1156.44 ;
     RECT  663.46 1204.96 683.14 1205.16 ;
     RECT  675.94 1319.2 683.14 1329.9 ;
     RECT  680.74 1288.54 683.62 1294.62 ;
     RECT  683.14 1319.2 683.62 1321.5 ;
     RECT  674.78 1189.84 685.06 1195.08 ;
     RECT  661.54 1412.02 685.06 1412.22 ;
     RECT  682.94 1258.72 685.34 1272.36 ;
     RECT  684.38 1295.26 686.02 1295.88 ;
     RECT  683.14 380.84 686.5 916.16 ;
     RECT  685.06 1189.84 686.5 1194.24 ;
     RECT  685.34 1253.68 686.5 1272.36 ;
     RECT  660.1 1367.5 686.98 1367.7 ;
     RECT  674.98 1228.48 687.46 1228.68 ;
     RECT  683.62 1321.3 687.94 1321.5 ;
     RECT  677.66 1423.78 687.94 1423.98 ;
     RECT  686.5 1257.88 688.7 1272.36 ;
     RECT  684.86 1209.16 688.9 1209.36 ;
     RECT  684.38 1330.12 688.9 1330.32 ;
     RECT  683.14 925.62 689.38 1156.44 ;
     RECT  689.38 925.62 689.86 1002.68 ;
     RECT  688.7 1357.84 691.1 1366.02 ;
     RECT  689.18 1245.28 691.58 1246.32 ;
     RECT  688.7 1296.1 692.06 1296.3 ;
     RECT  686.5 381.26 692.54 916.16 ;
     RECT  689.86 925.62 692.54 998.06 ;
     RECT  692.06 1296.1 693.98 1299.24 ;
     RECT  690.62 1397.32 694.18 1397.52 ;
     RECT  688.7 1257.88 695.14 1277.82 ;
     RECT  691.58 1416.22 695.14 1416.42 ;
     RECT  695.14 1257.88 696.1 1277.4 ;
     RECT  681.22 1449.32 696.38 1449.94 ;
     RECT  693.98 1296.1 696.86 1299.66 ;
     RECT  695.9 1383.04 697.34 1383.24 ;
     RECT  697.34 1201.18 697.82 1201.38 ;
     RECT  690.62 1231.42 698.3 1231.62 ;
     RECT  691.58 1241.5 698.3 1246.32 ;
     RECT  698.3 1231.42 699.26 1246.32 ;
     RECT  694.46 1337.26 699.26 1337.46 ;
     RECT  699.26 1336.84 699.74 1337.46 ;
     RECT  696.86 1296.1 700.22 1301.76 ;
     RECT  697.34 1383.04 700.9 1390.8 ;
     RECT  700.22 1296.1 701.86 1306.38 ;
     RECT  699.26 1223.86 702.62 1246.32 ;
     RECT  696.1 1257.88 702.62 1274.46 ;
     RECT  698.3 1322.56 702.62 1322.76 ;
     RECT  699.74 1333.9 702.62 1337.46 ;
     RECT  702.62 1322.56 702.82 1337.46 ;
     RECT  702.62 1223.86 704.26 1274.46 ;
     RECT  702.62 1401.52 704.26 1401.72 ;
     RECT  691.1 1355.74 705.02 1366.02 ;
     RECT  703.58 1283.92 706.46 1284.12 ;
     RECT  701.86 1296.1 706.46 1301.76 ;
     RECT  697.82 1193.62 707.42 1201.38 ;
     RECT  699.74 1210 707.42 1210.2 ;
     RECT  689.38 1012.98 708.58 1156.44 ;
     RECT  702.82 1330.12 709.34 1337.46 ;
     RECT  705.02 1351.96 709.34 1366.02 ;
     RECT  692.54 381.26 710.5 998.06 ;
     RECT  709.34 1330.12 710.5 1366.02 ;
     RECT  696.38 1448.56 711.26 1449.94 ;
     RECT  703.58 1315.42 711.94 1315.62 ;
     RECT  681.22 1459.4 713.18 1468.84 ;
     RECT  708.58 1033.56 713.38 1156.44 ;
     RECT  704.26 1223.86 713.66 1270.26 ;
     RECT  711.26 1447.3 713.66 1449.94 ;
     RECT  710.5 1330.12 713.86 1337.46 ;
     RECT  713.66 1446.46 713.86 1449.94 ;
     RECT  713.86 1330.12 714.82 1337.04 ;
     RECT  645 -70 715 178 ;
     RECT  677.86 1622 715 1870 ;
     RECT  713.66 1223.86 715.1 1274.46 ;
     RECT  706.46 1283.92 715.1 1301.76 ;
     RECT  698.78 1417.06 715.1 1417.26 ;
     RECT  700.9 1383.04 715.3 1383.24 ;
     RECT  715.1 1409.08 715.3 1417.26 ;
     RECT  714.82 1330.12 715.58 1330.32 ;
     RECT  715.1 1223.86 716.26 1301.76 ;
     RECT  713.38 1041.12 717.22 1156.44 ;
     RECT  710.5 1349.02 717.98 1366.02 ;
     RECT  717.98 1349.02 718.18 1374 ;
     RECT  716.26 1273.84 718.66 1301.76 ;
     RECT  672.38 220.82 719.19 221.02 ;
     RECT  588.81 255.26 719.19 255.46 ;
     RECT  588.81 269.96 719.19 270.16 ;
     RECT  658.46 327.5 719.19 356.26 ;
     RECT  710.5 381.26 719.19 990.5 ;
     RECT  588.81 1573.22 719.19 1579.3 ;
     RECT  713.86 1446.88 719.62 1449.94 ;
     RECT  707.42 1189.84 721.06 1210.2 ;
     RECT  718.66 1273.84 721.06 1278.24 ;
     RECT  721.06 1273.84 721.54 1276.98 ;
     RECT  713.18 1459.4 722.02 1469.76 ;
     RECT  713.66 1393.54 722.78 1393.74 ;
     RECT  718.18 1349.02 723.26 1358.04 ;
     RECT  719.19 215.36 723.46 990.5 ;
     RECT  723.46 215.36 724.81 916.58 ;
     RECT  719.19 1573.22 724.81 1583.92 ;
     RECT  712.7 1178.92 724.9 1179.12 ;
     RECT  723.46 926.46 725.18 990.5 ;
     RECT  715.58 1327.6 725.18 1330.32 ;
     RECT  717.22 1153.72 725.38 1156.44 ;
     RECT  722.78 1393.54 725.38 1397.94 ;
     RECT  725.18 926.46 725.86 995.12 ;
     RECT  723.26 1346.08 726.34 1358.04 ;
     RECT  715.3 1409.08 726.34 1410.96 ;
     RECT  708.58 1012.98 726.62 1021.58 ;
     RECT  719.62 1447.3 726.62 1449.94 ;
     RECT  722.02 1459.4 726.62 1468.84 ;
     RECT  724.81 381.26 726.82 916.58 ;
     RECT  718.18 1373.8 726.82 1374 ;
     RECT  725.18 1325.08 727.3 1330.32 ;
     RECT  726.34 1409.08 727.3 1409.28 ;
     RECT  716.26 1223.86 727.78 1263.96 ;
     RECT  726.62 1012.98 728.06 1023.26 ;
     RECT  726.34 1346.08 729.22 1356.36 ;
     RECT  726.62 1447.3 729.22 1468.84 ;
     RECT  725.38 1156.24 729.7 1156.44 ;
     RECT  727.3 1330.12 731.14 1330.32 ;
     RECT  729.22 1447.3 731.9 1449.94 ;
     RECT  727.78 1227.64 732.38 1263.96 ;
     RECT  718.66 1288.12 732.38 1301.76 ;
     RECT  732.38 1288.12 732.86 1302.18 ;
     RECT  715 0 733 178 ;
     RECT  715 1622 733 1800 ;
     RECT  725.86 932.76 733.34 995.12 ;
     RECT  732.86 1288.12 734.02 1306.38 ;
     RECT  733.34 932.76 734.3 1001.42 ;
     RECT  728.06 1010.46 734.3 1023.26 ;
     RECT  721.06 1189.84 734.3 1209.36 ;
     RECT  734.3 932.76 734.78 1023.26 ;
     RECT  732.38 1227.64 734.78 1266.06 ;
     RECT  721.54 1276.78 734.78 1276.98 ;
     RECT  717.22 1041.12 734.98 1145.06 ;
     RECT  734.78 1227.64 734.98 1276.98 ;
     RECT  729.22 1356.16 734.98 1356.36 ;
     RECT  734.3 1188.16 735.94 1209.78 ;
     RECT  734.98 1233.94 736.22 1276.98 ;
     RECT  734.02 1288.12 736.22 1302.18 ;
     RECT  734.78 932.76 736.42 1029.56 ;
     RECT  726.82 381.26 736.7 916.16 ;
     RECT  735.94 1188.58 736.7 1209.78 ;
     RECT  736.7 1188.58 737.38 1212.72 ;
     RECT  736.22 1233.94 737.86 1302.18 ;
     RECT  725.38 1397.74 737.86 1397.94 ;
     RECT  736.42 986.1 738.34 1029.56 ;
     RECT  737.86 1295.68 738.34 1302.18 ;
     RECT  731.9 1443.52 738.34 1449.94 ;
     RECT  737.38 1188.58 738.82 1195.08 ;
     RECT  729.22 1346.08 739.1 1346.28 ;
     RECT  725.66 1424.2 739.1 1424.4 ;
     RECT  737.86 1233.94 739.3 1281.6 ;
     RECT  731.42 1336.84 739.3 1337.04 ;
     RECT  739.1 1345.66 739.58 1346.28 ;
     RECT  739.58 1344.82 740.06 1346.28 ;
     RECT  738.34 986.94 740.54 1029.56 ;
     RECT  736.7 1171.36 740.54 1171.56 ;
     RECT  740.54 1412.86 741.5 1413.06 ;
     RECT  739.1 1424.2 741.5 1432.8 ;
     RECT  741.02 1368.34 742.18 1372.74 ;
     RECT  729.22 1459.4 742.94 1468.84 ;
     RECT  739.3 1274.26 743.62 1280.76 ;
     RECT  738.34 1299.88 744.38 1302.18 ;
     RECT  741.5 1412.86 744.38 1432.8 ;
     RECT  736.7 381.26 744.86 923.3 ;
     RECT  736.42 932.76 744.86 946.82 ;
     RECT  743.62 1274.26 745.06 1274.46 ;
     RECT  744.86 381.26 745.34 946.82 ;
     RECT  737.38 1209.16 745.54 1212.72 ;
     RECT  744.38 1299.88 746.02 1306.38 ;
     RECT  744.38 1408.66 746.02 1432.8 ;
     RECT  744.38 1390.6 746.3 1390.8 ;
     RECT  740.54 986.94 746.78 1031.66 ;
     RECT  745.54 1209.16 746.78 1209.36 ;
     RECT  740.06 1344.82 746.78 1349.22 ;
     RECT  746.02 1299.88 746.98 1302.18 ;
     RECT  746.78 1205.38 747.46 1209.36 ;
     RECT  742.18 1372.54 747.94 1372.74 ;
     RECT  746.78 986.94 748.7 1033.34 ;
     RECT  734.98 1042.38 748.7 1145.06 ;
     RECT  740.54 1171.36 749.38 1179.12 ;
     RECT  747.26 1299.46 749.66 1299.66 ;
     RECT  748.7 986.94 750.14 1145.06 ;
     RECT  742.94 1458.64 751.3 1468.84 ;
     RECT  741.5 1223.86 751.58 1224.06 ;
     RECT  739.3 1246.54 751.58 1261.44 ;
     RECT  750.14 1273.42 751.58 1273.62 ;
     RECT  746.78 1344.82 752.06 1356.78 ;
     RECT  738.34 1446.88 752.54 1449.94 ;
     RECT  745.34 381.26 752.74 947.24 ;
     RECT  752.06 1340.2 753.22 1356.78 ;
     RECT  752.74 925.16 753.5 947.24 ;
     RECT  736.42 955.86 753.5 976.64 ;
     RECT  752.54 1443.52 753.5 1449.94 ;
     RECT  753.5 925.16 753.98 976.64 ;
     RECT  750.14 985.68 753.98 1145.06 ;
     RECT  738.82 1194.88 753.98 1195.08 ;
     RECT  747.46 1205.38 753.98 1206 ;
     RECT  751.58 1223.86 754.66 1224.48 ;
     RECT  746.3 1390.6 754.66 1397.94 ;
     RECT  746.02 1408.66 755.14 1428.6 ;
     RECT  724.81 220.82 755.9 221.02 ;
     RECT  751.58 1246.54 756.1 1273.62 ;
     RECT  752.74 381.26 756.58 916.16 ;
     RECT  753.98 1189.84 756.58 1206 ;
     RECT  756.58 1189.84 756.86 1190.88 ;
     RECT  739.3 1233.94 756.86 1236.66 ;
     RECT  756.1 1246.54 756.86 1258.92 ;
     RECT  751.3 1459.4 757.34 1468.84 ;
     RECT  755.14 1408.66 757.54 1420.62 ;
     RECT  752.54 1329.7 757.82 1329.9 ;
     RECT  753.5 1443.1 758.3 1449.94 ;
     RECT  753.98 925.16 758.98 1145.06 ;
     RECT  753.22 1348.18 759.26 1356.78 ;
     RECT  757.54 1412.86 759.46 1420.62 ;
     RECT  754.66 1224.28 760.22 1224.48 ;
     RECT  756.86 1233.94 760.22 1258.92 ;
     RECT  758.98 925.16 760.42 1144.22 ;
     RECT  749.66 1294.84 761.18 1299.66 ;
     RECT  749.38 1171.36 761.38 1171.56 ;
     RECT  761.18 1288.12 761.38 1299.66 ;
     RECT  759.26 1348.18 761.38 1361.32 ;
     RECT  758.78 1310.38 762.82 1310.58 ;
     RECT  754.66 1390.6 762.82 1390.8 ;
     RECT  760.42 925.16 763.3 1143.38 ;
     RECT  756.86 1186.48 764.26 1190.88 ;
     RECT  758.3 1435.54 764.26 1449.94 ;
     RECT  764.26 1435.54 764.54 1447.5 ;
     RECT  756.58 1205.8 765.02 1206 ;
     RECT  763.3 946.62 766.18 1143.38 ;
     RECT  760.22 1224.28 766.18 1258.92 ;
     RECT  756.1 1269.64 766.18 1273.62 ;
     RECT  759.46 1412.86 766.18 1413.06 ;
     RECT  762.62 1378.84 766.46 1379.04 ;
     RECT  757.34 1459.4 767.14 1473.54 ;
     RECT  766.46 1375.06 767.9 1379.04 ;
     RECT  764.26 1186.48 769.06 1186.68 ;
     RECT  756.58 381.26 769.82 592.72 ;
     RECT  756.58 601.34 769.82 916.16 ;
     RECT  765.02 1202.02 769.82 1206 ;
     RECT  766.18 1224.28 769.82 1231.62 ;
     RECT  768.86 1318.36 769.82 1318.56 ;
     RECT  757.82 1329.7 769.82 1330.66 ;
     RECT  766.18 1246.96 770.3 1258.92 ;
     RECT  766.18 946.62 770.5 1137.5 ;
     RECT  761.38 1299.46 770.98 1299.66 ;
     RECT  769.82 1201.18 771.46 1206 ;
     RECT  769.82 1221.76 771.46 1231.62 ;
     RECT  764.06 1340.96 771.74 1341.16 ;
     RECT  766.18 1273.42 772.42 1273.62 ;
     RECT  769.82 1318.36 772.9 1330.66 ;
     RECT  764.54 1432.18 773.18 1447.5 ;
     RECT  767.14 1459.4 773.18 1468.84 ;
     RECT  772.9 1329.7 773.38 1330.66 ;
     RECT  770.5 946.62 774.34 1137.46 ;
     RECT  771.46 1224.28 775.3 1231.62 ;
     RECT  770.3 1246.96 775.3 1262.28 ;
     RECT  768.86 1416.64 777.02 1416.84 ;
     RECT  773.18 1432.18 777.22 1468.84 ;
     RECT  767.9 1371.28 777.5 1379.04 ;
     RECT  777.5 1371.28 777.7 1382.82 ;
     RECT  777.22 1446.88 777.7 1468.84 ;
     RECT  772.9 1318.36 778.66 1319.32 ;
     RECT  769.82 381.26 779.42 916.16 ;
     RECT  763.3 925.16 779.42 934.64 ;
     RECT  771.74 1340.96 779.42 1345.44 ;
     RECT  761.38 1356.58 779.42 1361.32 ;
     RECT  775.3 1224.28 779.62 1224.48 ;
     RECT  774.34 1133.1 780.86 1137.46 ;
     RECT  779.42 381.26 781.54 934.64 ;
     RECT  774.34 946.62 781.82 1124.06 ;
     RECT  779.42 1340.96 782.02 1361.32 ;
     RECT  777.02 1412.86 782.02 1416.84 ;
     RECT  777.22 1432.18 782.5 1435.74 ;
     RECT  774.62 1304.5 782.78 1305.12 ;
     RECT  777.7 1379.26 782.78 1382.82 ;
     RECT  782.78 1379.26 782.98 1384.08 ;
     RECT  782.02 1416.64 783.94 1416.84 ;
     RECT  782.5 1435.54 784.9 1435.74 ;
     RECT  761.38 1288.12 785.18 1288.32 ;
     RECT  782.78 1296.94 785.18 1305.12 ;
     RECT  785.18 1288.12 786.34 1305.12 ;
     RECT  777.7 1454.86 786.34 1468.84 ;
     RECT  786.34 1300.72 786.82 1305.12 ;
     RECT  755.9 220.82 787.19 221.86 ;
     RECT  724.81 255.26 787.19 255.46 ;
     RECT  724.81 269.96 787.19 270.16 ;
     RECT  786.62 284.24 787.19 284.44 ;
     RECT  724.81 327.5 787.19 356.26 ;
     RECT  746.78 370.76 787.19 370.96 ;
     RECT  781.54 381.26 787.19 916.16 ;
     RECT  724.81 1573.22 787.19 1579.3 ;
     RECT  773.38 1330.46 788.06 1330.66 ;
     RECT  782.98 1379.26 788.26 1382.82 ;
     RECT  786.62 1278.46 788.74 1278.66 ;
     RECT  781.82 944.9 789.5 1124.06 ;
     RECT  780.86 1133.1 789.5 1141.66 ;
     RECT  775.3 1249.9 789.5 1262.28 ;
     RECT  789.5 1248.22 789.7 1269.84 ;
     RECT  789.7 1257.88 790.66 1258.5 ;
     RECT  787.19 219.14 791.9 916.16 ;
     RECT  781.54 925.16 791.9 934.64 ;
     RECT  788.06 1330.46 791.9 1331.16 ;
     RECT  791.9 219.14 792.81 934.64 ;
     RECT  787.19 1573.22 792.81 1580.14 ;
     RECT  792.81 601.34 793.82 934.64 ;
     RECT  791.9 1330.04 793.82 1331.16 ;
     RECT  782.02 1340.96 793.82 1351.74 ;
     RECT  793.82 1330.04 795.46 1351.74 ;
     RECT  790.94 1405.3 796.22 1405.5 ;
     RECT  789.7 1269.64 797.18 1269.84 ;
     RECT  790.46 1280.98 797.18 1281.18 ;
     RECT  789.98 1378.84 797.18 1379.04 ;
     RECT  796.22 1405.3 797.18 1409.7 ;
     RECT  794.3 1233.1 797.38 1239.6 ;
     RECT  795.46 1340.96 797.38 1349.64 ;
     RECT  796.7 1189.84 798.14 1190.04 ;
     RECT  789.5 1198.66 798.14 1198.86 ;
     RECT  797.38 1239.4 798.14 1239.6 ;
     RECT  789.7 1248.22 798.14 1248.42 ;
     RECT  786.82 1300.72 798.14 1304.28 ;
     RECT  787.1 1440.16 798.14 1443.3 ;
     RECT  797.18 1377.16 798.34 1379.04 ;
     RECT  798.14 1440.16 798.34 1447.5 ;
     RECT  793.82 601.34 799.1 935.06 ;
     RECT  789.5 944.9 799.1 1141.66 ;
     RECT  797.18 1400.26 799.1 1409.7 ;
     RECT  791.42 1424.2 799.1 1424.4 ;
     RECT  795.26 1220.5 800.06 1220.7 ;
     RECT  800.06 1220.5 800.26 1228.26 ;
     RECT  790.66 1258.3 800.26 1258.5 ;
     RECT  798.14 1189.84 800.74 1198.86 ;
     RECT  799.1 1400.26 801.5 1410.12 ;
     RECT  797.18 1269.64 802.94 1281.18 ;
     RECT  733 -70 803 178 ;
     RECT  733 1622 803 1870 ;
     RECT  802.94 1265.44 804.38 1281.18 ;
     RECT  799.1 601.34 804.58 1141.66 ;
     RECT  804.58 601.34 805.06 1127.8 ;
     RECT  795.46 1330.04 805.06 1331.16 ;
     RECT  798.34 1378.84 805.34 1379.04 ;
     RECT  805.06 601.34 805.54 1034.18 ;
     RECT  798.14 1299.88 806.78 1304.28 ;
     RECT  804.38 1265.44 806.98 1287.48 ;
     RECT  805.54 601.34 807.46 1032.5 ;
     RECT  800.26 1227.64 807.46 1228.26 ;
     RECT  806.78 1296.52 807.74 1304.28 ;
     RECT  805.34 1378.84 807.94 1382.82 ;
     RECT  806.98 1265.44 808.42 1284.54 ;
     RECT  807.94 1378.84 808.42 1379.04 ;
     RECT  778.66 1319.12 808.7 1319.32 ;
     RECT  805.06 1043.64 809.38 1127.8 ;
     RECT  797.38 1340.96 809.66 1348.8 ;
     RECT  792.81 381.26 809.86 592.72 ;
     RECT  809.38 1076.4 809.86 1127.8 ;
     RECT  807.46 1228.06 810.14 1228.26 ;
     RECT  798.14 1239.4 810.14 1248.42 ;
     RECT  798.34 1442.68 810.34 1447.5 ;
     RECT  801.5 1400.26 811.1 1410.54 ;
     RECT  799.1 1424.2 811.1 1425.66 ;
     RECT  811.1 1400.26 811.3 1425.66 ;
     RECT  805.34 1208.74 812.54 1208.94 ;
     RECT  810.34 1443.1 812.74 1447.5 ;
     RECT  808.7 1314.58 813.5 1319.32 ;
     RECT  805.06 1330.04 813.5 1330.24 ;
     RECT  810.14 1228.06 813.98 1248.42 ;
     RECT  807.74 1296.52 813.98 1304.7 ;
     RECT  813.5 1314.58 813.98 1330.24 ;
     RECT  809.86 1078.08 815.14 1127.8 ;
     RECT  800.74 1193.62 815.14 1198.86 ;
     RECT  809.66 1340.96 815.14 1352.58 ;
     RECT  808.7 1182.7 815.9 1182.9 ;
     RECT  815.14 1197.4 815.9 1198.86 ;
     RECT  812.54 1208.74 815.9 1212.72 ;
     RECT  815.14 1078.08 816.1 1110.2 ;
     RECT  815.14 1122.6 816.58 1127.8 ;
     RECT  811.3 1400.26 816.58 1416.84 ;
     RECT  809.86 404.78 816.86 592.72 ;
     RECT  807.46 601.34 816.86 1027.04 ;
     RECT  813.98 1296.52 816.86 1330.24 ;
     RECT  815.14 1340.96 816.86 1348.8 ;
     RECT  808.42 1265.44 817.06 1281.18 ;
     RECT  817.06 1265.44 817.54 1265.64 ;
     RECT  817.06 1277.2 818.3 1281.18 ;
     RECT  816.86 1296.52 818.3 1348.8 ;
     RECT  818.3 1277.2 818.5 1348.8 ;
     RECT  816.1 1095.72 818.98 1110.2 ;
     RECT  809.38 1043.64 819.26 1063.58 ;
     RECT  815.9 1182.7 819.26 1184.5 ;
     RECT  816.1 1078.08 819.46 1087.1 ;
     RECT  812.74 1443.1 819.46 1447.08 ;
     RECT  818.98 1095.72 819.94 1097.6 ;
     RECT  817.82 1382.2 820.42 1386.6 ;
     RECT  818.98 1106.22 820.9 1110.2 ;
     RECT  803 0 821 178 ;
     RECT  803 1622 821 1800 ;
     RECT  816.86 404.78 821.38 1027.04 ;
     RECT  818.5 1277.2 821.38 1319.32 ;
     RECT  819.94 1095.72 821.86 1096.76 ;
     RECT  816.86 1371.28 821.86 1371.48 ;
     RECT  813.98 1228.06 822.14 1250.94 ;
     RECT  819.46 1081.86 822.34 1087.1 ;
     RECT  821.86 1095.72 823.3 1096.34 ;
     RECT  820.9 1108.32 823.3 1108.52 ;
     RECT  819.26 1040.66 824.06 1063.58 ;
     RECT  823.3 1096.14 824.26 1096.34 ;
     RECT  820.42 1386.4 824.74 1386.6 ;
     RECT  786.34 1459.4 824.74 1468.84 ;
     RECT  822.14 1224.28 825.22 1250.94 ;
     RECT  821.38 404.78 825.7 982.48 ;
     RECT  819.26 1182.28 825.98 1184.5 ;
     RECT  821.38 1277.2 826.18 1309.74 ;
     RECT  811.3 1425.46 827.14 1425.66 ;
     RECT  815.9 1197.4 827.42 1212.72 ;
     RECT  825.98 1176.82 828.1 1184.5 ;
     RECT  825.5 1266.28 828.38 1266.48 ;
     RECT  816.58 1400.26 829.34 1416.42 ;
     RECT  826.18 1277.2 829.54 1278.66 ;
     RECT  827.42 1197.4 830.02 1213.48 ;
     RECT  828.38 1262.5 830.02 1266.48 ;
     RECT  821.38 991.94 831.26 1027.04 ;
     RECT  824.06 1040.24 831.26 1063.58 ;
     RECT  821.38 1319.12 831.26 1319.32 ;
     RECT  818.5 1330.04 831.26 1348.8 ;
     RECT  825.7 601.34 831.74 982.48 ;
     RECT  831.26 1319.12 831.94 1348.8 ;
     RECT  829.54 1278.46 832.42 1278.66 ;
     RECT  830.02 1202.86 832.9 1213.48 ;
     RECT  829.34 1400.26 833.38 1418.1 ;
     RECT  819.46 1443.1 834.14 1446.24 ;
     RECT  792.81 327.5 834.62 356.26 ;
     RECT  792.81 370.76 834.62 370.96 ;
     RECT  831.94 1319.12 834.82 1345.02 ;
     RECT  830.02 1262.5 835.78 1262.7 ;
     RECT  826.18 1289.3 835.78 1309.74 ;
     RECT  833.38 1417.9 835.78 1418.1 ;
     RECT  825.22 1234.28 836.54 1250.94 ;
     RECT  834.14 1439.32 836.74 1447.08 ;
     RECT  828.1 1182.28 837.22 1184.5 ;
     RECT  836.74 1446.88 838.18 1447.08 ;
     RECT  831.74 601.34 839.42 983.36 ;
     RECT  831.26 991.94 839.42 1063.58 ;
     RECT  835.78 1289.3 839.62 1306.8 ;
     RECT  839.62 1289.3 839.9 1304.7 ;
     RECT  839.9 1281.82 840.1 1304.7 ;
     RECT  837.22 1183.88 840.86 1184.5 ;
     RECT  825.7 404.78 842.02 592.72 ;
     RECT  834.82 1319.12 842.02 1343.26 ;
     RECT  839.9 1381.36 842.02 1381.56 ;
     RECT  840.38 1194.88 842.78 1195.08 ;
     RECT  832.9 1204.54 842.78 1213.48 ;
     RECT  833.38 1400.26 842.78 1405.92 ;
     RECT  792.81 220.82 843.74 221.86 ;
     RECT  842.78 1194.88 844.22 1213.48 ;
     RECT  809.86 381.26 844.9 395.74 ;
     RECT  825.22 1224.28 845.18 1224.48 ;
     RECT  836.54 1234.28 845.18 1254.72 ;
     RECT  840.86 1431.76 845.18 1431.96 ;
     RECT  842.02 1319.12 845.66 1319.32 ;
     RECT  792.81 1573.22 845.86 1579.3 ;
     RECT  845.18 1224.28 846.14 1254.72 ;
     RECT  844.22 1265.44 846.14 1265.64 ;
     RECT  842.78 1390.18 846.14 1405.92 ;
     RECT  843.26 1420.42 846.14 1420.62 ;
     RECT  845.18 1431.34 846.14 1431.96 ;
     RECT  839.42 601.34 846.34 1063.58 ;
     RECT  844.22 1194.88 846.62 1215.58 ;
     RECT  846.14 1224.28 846.62 1265.64 ;
     RECT  840.1 1281.82 846.62 1296.3 ;
     RECT  846.14 1420.42 847.3 1431.96 ;
     RECT  846.62 1194.88 848.06 1265.64 ;
     RECT  846.62 1277.62 848.06 1296.3 ;
     RECT  843.26 1447.3 848.06 1447.5 ;
     RECT  843.26 1375.48 848.74 1375.68 ;
     RECT  847.3 1424.2 848.74 1431.96 ;
     RECT  848.06 1194.88 849.02 1296.3 ;
     RECT  822.34 1084.38 849.5 1087.1 ;
     RECT  846.34 601.34 849.7 994.7 ;
     RECT  849.02 1194.88 849.7 1300.08 ;
     RECT  849.7 1273 850.46 1300.08 ;
     RECT  850.46 1273 850.66 1303.44 ;
     RECT  842.02 404.78 850.94 587.26 ;
     RECT  845.86 1574.06 850.94 1579.3 ;
     RECT  849.5 1084.38 851.14 1087.9 ;
     RECT  846.14 1390.18 851.62 1408.44 ;
     RECT  840.86 1183.88 851.9 1185.34 ;
     RECT  849.7 1194.88 851.9 1261.86 ;
     RECT  842.02 1330.04 852.1 1343.26 ;
     RECT  850.66 1277.62 852.58 1303.44 ;
     RECT  851.62 1390.18 852.58 1405.92 ;
     RECT  848.74 1424.2 853.06 1425.24 ;
     RECT  851.14 1086.9 853.34 1087.9 ;
     RECT  849.7 601.34 854.02 992.56 ;
     RECT  850.94 1574.06 854.02 1583.08 ;
     RECT  846.34 1003.7 854.98 1063.58 ;
     RECT  852.58 1277.62 854.98 1282.02 ;
     RECT  852.58 1393.96 854.98 1405.92 ;
     RECT  854.02 601.34 855.46 982.48 ;
     RECT  854.98 1401.94 855.46 1405.92 ;
     RECT  853.06 1425.04 855.46 1425.24 ;
     RECT  848.06 1443.1 855.94 1447.5 ;
     RECT  854.98 1003.7 856.42 1049.72 ;
     RECT  854.78 1173.8 856.42 1174 ;
     RECT  851.9 1183.88 857.38 1261.86 ;
     RECT  854.98 1277.62 857.38 1277.82 ;
     RECT  855.94 1443.1 857.38 1443.3 ;
     RECT  855.46 602.6 858.34 982.48 ;
     RECT  853.34 1086.9 858.34 1090.84 ;
     RECT  852.1 1330.04 858.34 1342.42 ;
     RECT  845.66 1314.58 858.62 1319.32 ;
     RECT  850.94 404.78 859.3 588.52 ;
     RECT  856.42 1003.7 860.26 1028.72 ;
     RECT  292.22 1529.96 860.26 1551.58 ;
     RECT  857.38 1261.66 861.5 1261.86 ;
     RECT  854.98 1061.66 861.7 1063.58 ;
     RECT  857.38 1183.88 861.7 1250.94 ;
     RECT  858.34 934.44 862.18 982.48 ;
     RECT  856.42 1039.82 863.14 1049.72 ;
     RECT  855.46 1401.94 863.14 1402.14 ;
     RECT  860.26 1003.7 865.54 1026.58 ;
     RECT  854.02 1574.06 865.82 1580.98 ;
     RECT  844.9 382.94 866.02 395.74 ;
     RECT  865.54 1003.7 866.02 1006.04 ;
     RECT  852.58 1291.82 866.78 1303.44 ;
     RECT  861.7 1183.88 867.74 1247.16 ;
     RECT  858.34 602.6 870.82 925.78 ;
     RECT  866.02 382.94 871.3 394.9 ;
     RECT  866.78 1284.34 871.3 1303.44 ;
     RECT  867.74 1182.62 871.78 1247.16 ;
     RECT  858.34 1342.22 872.54 1342.42 ;
     RECT  862.18 934.44 873.22 978.28 ;
     RECT  871.3 1284.34 873.98 1303.36 ;
     RECT  861.5 1261.66 874.18 1266.06 ;
     RECT  280.22 1486.7 874.66 1515.88 ;
     RECT  865.82 1574.06 874.66 1583.08 ;
     RECT  873.98 1281.32 874.94 1303.36 ;
     RECT  873.22 939.02 875.42 978.28 ;
     RECT  854.02 991.52 875.42 992.56 ;
     RECT  872.54 1342.22 875.62 1345.44 ;
     RECT  792.81 255.26 875.9 255.46 ;
     RECT  792.81 269.96 875.9 270.16 ;
     RECT  871.3 382.94 876.1 388.18 ;
     RECT  874.18 1261.66 876.86 1261.86 ;
     RECT  875.42 939.02 877.06 992.56 ;
     RECT  868.7 1420.42 877.06 1420.62 ;
     RECT  874.94 1274.6 880.9 1303.36 ;
     RECT  865.54 1016.3 881.18 1026.58 ;
     RECT  870.82 602.6 881.66 899.32 ;
     RECT  870.82 909.62 881.66 925.78 ;
     RECT  877.06 939.02 881.66 992.14 ;
     RECT  866.02 1003.7 882.14 1005.16 ;
     RECT  881.18 1015.04 882.14 1026.58 ;
     RECT  871.78 1220.42 882.14 1247.16 ;
     RECT  876.86 1256.12 882.14 1261.86 ;
     RECT  858.62 1314.16 882.14 1319.32 ;
     RECT  859.3 404.78 882.34 587.26 ;
     RECT  748.7 1601.78 882.34 1601.98 ;
     RECT  804.58 1137.26 882.62 1141.66 ;
     RECT  882.62 1137.26 884.54 1150.06 ;
     RECT  881.66 909.62 885.5 992.14 ;
     RECT  885.5 908.36 887.42 992.14 ;
     RECT  882.14 1220.42 887.42 1261.86 ;
     RECT  880.9 1274.6 887.42 1281.52 ;
     RECT  880.9 1291.82 887.9 1303.36 ;
     RECT  882.14 1312.82 887.9 1319.32 ;
     RECT  882.34 583.7 888.38 587.26 ;
     RECT  881.66 602.18 888.38 899.32 ;
     RECT  888.38 583.7 888.58 899.32 ;
     RECT  875.62 1342.22 888.86 1342.42 ;
     RECT  860.26 1529.96 889.54 1544.44 ;
     RECT  887.42 908.36 890.3 995.08 ;
     RECT  882.14 1003.7 890.3 1026.58 ;
     RECT  874.66 1486.7 890.5 1515.46 ;
     RECT  821 -70 891 178 ;
     RECT  821 1622 891 1870 ;
     RECT  863.14 1039.82 891.26 1048 ;
     RECT  861.7 1061.66 891.26 1061.86 ;
     RECT  890.5 1500.98 891.46 1515.46 ;
     RECT  888.58 583.7 891.94 584.32 ;
     RECT  858.34 1330.04 892.7 1332.76 ;
     RECT  888.86 1342.22 892.7 1342.84 ;
     RECT  892.7 1330.04 892.9 1342.84 ;
     RECT  891.26 1039.82 893.18 1061.86 ;
     RECT  888.58 595.46 895.3 899.32 ;
     RECT  898.94 1173.38 899.42 1173.58 ;
     RECT  871.78 1182.62 899.42 1210.96 ;
     RECT  899.42 1173.38 899.9 1210.96 ;
     RECT  899.9 1170.02 900.86 1210.96 ;
     RECT  824.74 1459.4 901.035 1459.6 ;
     RECT  824.74 1468.64 901.035 1468.84 ;
     RECT  890.5 1486.7 901.035 1487.32 ;
     RECT  891.46 1500.98 901.035 1508.32 ;
     RECT  889.54 1529.96 901.035 1537.3 ;
     RECT  874.66 1574.06 901.035 1580.98 ;
     RECT  884.54 1137.26 902.3 1155.52 ;
     RECT  900.86 1166.24 902.78 1210.96 ;
     RECT  887.42 1220.42 902.78 1281.52 ;
     RECT  901.035 1372.04 902.965 1583.92 ;
     RECT  858.34 1090.64 903.46 1090.84 ;
     RECT  902.3 1137.26 903.74 1155.94 ;
     RECT  902.78 1166.24 903.74 1281.52 ;
     RECT  902.965 1529.96 903.94 1531 ;
     RECT  903.74 1137.26 904.22 1281.52 ;
     RECT  904.22 1136.84 904.7 1281.52 ;
     RECT  887.9 1291.82 904.7 1319.32 ;
     RECT  892.9 1330.46 904.7 1342.84 ;
     RECT  890.3 908.36 904.9 1026.58 ;
     RECT  904.9 908.36 906.14 1024.9 ;
     RECT  902.965 1459.4 906.34 1459.6 ;
     RECT  895.3 602.6 906.62 899.32 ;
     RECT  906.14 907.94 906.62 1024.9 ;
     RECT  816.58 1127.6 907.1 1127.8 ;
     RECT  904.7 1291.82 907.3 1342.84 ;
     RECT  893.18 1039.82 907.58 1063.54 ;
     RECT  907.1 1125.08 907.58 1127.8 ;
     RECT  904.7 1136.42 907.58 1281.52 ;
     RECT  882.34 404.78 907.78 574.24 ;
     RECT  902.965 1492.58 907.78 1493.62 ;
     RECT  899.42 1107.02 908.06 1107.22 ;
     RECT  907.58 1125.08 908.06 1281.52 ;
     RECT  908.06 1125.08 908.26 1282.36 ;
     RECT  907.3 1301.06 908.26 1342.84 ;
     RECT  908.26 1125.08 908.54 1215.58 ;
     RECT  782.02 1361.12 908.54 1361.32 ;
     RECT  891 0 909 178 ;
     RECT  891 1622 909 1800 ;
     RECT  906.62 602.6 909.02 1024.9 ;
     RECT  908.54 1124.24 909.02 1215.58 ;
     RECT  907.78 1493.42 909.7 1493.62 ;
     RECT  907.58 1037.3 909.98 1063.54 ;
     RECT  908.54 1361.12 909.98 1363 ;
     RECT  909.98 1037.3 910.46 1068.16 ;
     RECT  908.26 1224.62 910.46 1282.36 ;
     RECT  907.3 1291.82 910.46 1292.02 ;
     RECT  902.965 1519.04 911.42 1519.24 ;
     RECT  902.965 1468.64 912.86 1468.84 ;
     RECT  909.02 595.04 913.34 1024.9 ;
     RECT  908.06 1107.02 913.34 1108.9 ;
     RECT  909.02 1121.3 913.34 1215.58 ;
     RECT  902.965 1377.92 913.82 1378.12 ;
     RECT  903.94 1530.8 913.82 1531 ;
     RECT  908.26 1325 914.3 1342.84 ;
     RECT  909.98 1352.72 914.3 1363 ;
     RECT  913.82 1377.92 914.3 1385.68 ;
     RECT  912.86 1466.12 915.74 1468.84 ;
     RECT  910.46 1037.3 916.22 1073.2 ;
     RECT  915.74 1455.62 916.42 1468.84 ;
     RECT  913.34 595.04 916.7 1026.16 ;
     RECT  916.22 1036.88 916.7 1073.2 ;
     RECT  913.34 1107.02 916.7 1215.58 ;
     RECT  891.94 584.12 917.18 584.32 ;
     RECT  916.7 595.04 917.18 1073.2 ;
     RECT  914.3 1325 917.18 1363 ;
     RECT  914.3 1377.08 917.18 1385.68 ;
     RECT  911.42 1519.04 917.86 1520.08 ;
     RECT  917.18 1325 918.14 1385.68 ;
     RECT  913.82 1530.8 918.62 1534.36 ;
     RECT  915.74 1422.02 918.82 1422.22 ;
     RECT  916.7 1097.78 919.1 1215.58 ;
     RECT  910.46 1224.62 919.1 1292.02 ;
     RECT  908.26 1301.06 919.1 1313.02 ;
     RECT  917.18 1553.06 919.1 1553.26 ;
     RECT  917.18 584.12 919.58 1073.2 ;
     RECT  919.1 1224.2 919.58 1313.02 ;
     RECT  918.14 1325 919.58 1386.1 ;
     RECT  919.1 1093.16 920.54 1215.58 ;
     RECT  919.58 1224.2 920.54 1386.1 ;
     RECT  917.86 1519.46 920.74 1520.08 ;
     RECT  920.54 1093.16 921.02 1386.1 ;
     RECT  918.62 1530.8 921.22 1539.4 ;
     RECT  921.02 1090.64 921.5 1386.1 ;
     RECT  916.42 1467.38 921.98 1468.84 ;
     RECT  921.22 1531.22 921.98 1539.4 ;
     RECT  919.1 1550.54 921.98 1554.52 ;
     RECT  909 -70 922.46 178 ;
     RECT  843.74 216.2 923.19 221.86 ;
     RECT  875.9 255.26 923.19 270.16 ;
     RECT  792.81 284.24 923.19 284.44 ;
     RECT  834.62 327.5 923.19 370.96 ;
     RECT  876.1 383.36 923.19 388.18 ;
     RECT  907.78 406.46 923.19 574.24 ;
     RECT  919.58 584.12 923.19 1073.62 ;
     RECT  921.5 1084.76 923.19 1386.1 ;
     RECT  902.965 1574.06 923.19 1580.98 ;
     RECT  921.98 1531.22 924.1 1554.52 ;
     RECT  924.1 1535 924.58 1554.52 ;
     RECT  909 1622 924.86 1870 ;
     RECT  916.42 1455.62 925.82 1455.82 ;
     RECT  920.74 1519.46 926.02 1519.66 ;
     RECT  924.58 1535 926.02 1554.1 ;
     RECT  923.42 1435.04 926.3 1435.24 ;
     RECT  925.82 1452.68 926.3 1455.82 ;
     RECT  921.98 1467.38 926.3 1475.14 ;
     RECT  921.02 1485.02 926.3 1486.9 ;
     RECT  926.3 1448.06 926.78 1455.82 ;
     RECT  926.3 1467.38 926.78 1486.9 ;
     RECT  925.82 1410.26 928.7 1410.46 ;
     RECT  923.19 215.36 928.81 1386.1 ;
     RECT  923.19 1574.06 928.81 1583.92 ;
     RECT  926.3 1429.58 929.66 1435.24 ;
     RECT  926.78 1448.06 929.66 1486.9 ;
     RECT  928.81 1090.64 929.86 1287.4 ;
     RECT  929.66 1424.54 929.86 1486.9 ;
     RECT  929.86 1236.38 930.34 1287.4 ;
     RECT  928.81 599.24 930.82 1072.78 ;
     RECT  930.34 1236.38 930.82 1283.62 ;
     RECT  928.7 1410.26 931.1 1410.88 ;
     RECT  930.82 1236.38 931.78 1240.78 ;
     RECT  930.82 613.94 932.26 1072.78 ;
     RECT  928.81 1296.44 932.54 1386.1 ;
     RECT  932.26 614.78 932.74 1072.78 ;
     RECT  932.54 1296.44 933.22 1388.2 ;
     RECT  929.86 1424.54 933.7 1458.76 ;
     RECT  926.02 1535 933.7 1550.74 ;
     RECT  931.1 1410.26 933.98 1414.66 ;
     RECT  933.7 1424.54 933.98 1457.92 ;
     RECT  930.82 599.24 935.14 604.48 ;
     RECT  933.7 1546.34 935.14 1550.74 ;
     RECT  935.14 1550.54 935.42 1550.74 ;
     RECT  933.98 1561.46 935.42 1561.66 ;
     RECT  930.82 1249.4 935.62 1283.62 ;
     RECT  933.98 1410.26 935.62 1457.92 ;
     RECT  932.06 1399.76 935.9 1399.96 ;
     RECT  935.62 1410.26 935.9 1452.88 ;
     RECT  933.7 1535 936.38 1535.2 ;
     RECT  936.38 1531.22 936.58 1535.2 ;
     RECT  932.74 916.76 937.54 1072.78 ;
     RECT  933.22 1296.44 937.54 1318.48 ;
     RECT  937.54 1296.44 937.82 1300.42 ;
     RECT  937.54 1309.04 938.02 1318.48 ;
     RECT  929.86 1467.38 938.02 1486.9 ;
     RECT  935.9 1399.76 938.5 1452.88 ;
     RECT  936.58 1531.22 939.46 1534.78 ;
     RECT  935.42 1550.54 939.46 1561.66 ;
     RECT  929.86 1090.64 940.22 1227.34 ;
     RECT  937.54 916.76 940.42 950.56 ;
     RECT  937.54 959.6 940.7 1072.78 ;
     RECT  940.22 1083.92 940.7 1227.34 ;
     RECT  913.34 1508.96 940.7 1509.16 ;
     RECT  932.74 614.78 942.62 907.72 ;
     RECT  940.7 959.6 942.82 1227.34 ;
     RECT  935.14 602.6 943.1 604.48 ;
     RECT  942.62 614.78 943.1 908.14 ;
     RECT  931.78 1238.06 943.1 1240.78 ;
     RECT  938.02 1474.52 943.58 1486.9 ;
     RECT  927.74 1497.2 943.58 1497.4 ;
     RECT  943.1 602.6 943.78 908.14 ;
     RECT  928.81 406.46 944.26 584.74 ;
     RECT  939.46 1554.32 945.22 1561.66 ;
     RECT  943.1 1237.22 945.98 1240.78 ;
     RECT  935.62 1251.5 945.98 1283.62 ;
     RECT  942.82 1032.68 946.66 1227.34 ;
     RECT  945.98 1237.22 947.14 1283.62 ;
     RECT  938.5 1399.76 947.14 1441.12 ;
     RECT  943.78 615.62 947.9 908.14 ;
     RECT  933.22 1327.52 947.9 1388.2 ;
     RECT  947.14 1399.76 947.9 1399.96 ;
     RECT  943.58 1474.52 947.9 1497.4 ;
     RECT  947.14 1237.22 948.1 1255.9 ;
     RECT  947.14 1271.66 948.1 1283.62 ;
     RECT  940.42 918.02 948.38 950.56 ;
     RECT  942.82 959.6 948.38 1023.64 ;
     RECT  948.1 1272.5 948.86 1283.62 ;
     RECT  937.82 1295.6 948.86 1300.42 ;
     RECT  946.66 1078.46 949.06 1227.34 ;
     RECT  948.38 918.02 949.54 1023.64 ;
     RECT  949.06 1078.46 950.02 1200.88 ;
     RECT  945.22 1561.46 950.02 1561.66 ;
     RECT  939.46 1534.58 950.5 1534.78 ;
     RECT  950.02 1078.46 950.98 1198.78 ;
     RECT  944.26 583.7 951.94 584.74 ;
     RECT  947.14 1410.68 951.94 1441.12 ;
     RECT  947.9 1466.96 951.94 1497.4 ;
     RECT  951.94 1474.52 952.42 1497.4 ;
     RECT  947.9 615.62 953.66 908.56 ;
     RECT  949.54 918.02 953.66 928.3 ;
     RECT  938.5 1452.68 954.62 1452.88 ;
     RECT  952.42 1474.52 954.82 1490.68 ;
     RECT  949.06 1211.18 955.1 1227.34 ;
     RECT  946.66 1032.68 955.58 1069 ;
     RECT  950.98 1078.46 955.58 1084.54 ;
     RECT  948.1 1240.58 955.58 1255.9 ;
     RECT  938.02 1312.82 955.58 1318.48 ;
     RECT  947.9 1327.52 955.58 1399.96 ;
     RECT  950.98 1093.16 956.26 1198.78 ;
     RECT  940.7 1508.54 957.02 1509.16 ;
     RECT  954.62 1451.84 957.22 1452.88 ;
     RECT  956.26 1093.16 957.7 1113.52 ;
     RECT  955.1 1211.18 957.7 1230.7 ;
     RECT  943.78 602.6 957.98 606.58 ;
     RECT  953.66 615.62 957.98 928.3 ;
     RECT  954.82 1477.04 958.18 1490.68 ;
     RECT  955.58 1032.68 958.46 1084.54 ;
     RECT  957.7 1211.18 958.66 1227.34 ;
     RECT  951.94 1413.62 958.66 1441.12 ;
     RECT  957.98 602.6 958.94 928.3 ;
     RECT  949.54 939.44 958.94 1023.64 ;
     RECT  958.46 1032.26 958.94 1084.54 ;
     RECT  958.66 1413.62 959.14 1440.7 ;
     RECT  951.94 584.54 960.38 584.74 ;
     RECT  958.18 1477.04 960.58 1490.26 ;
     RECT  948.86 1272.5 960.86 1300.42 ;
     RECT  957.7 1093.16 961.54 1113.1 ;
     RECT  955.58 1240.58 962.3 1259.26 ;
     RECT  960.86 1463.6 963.26 1463.8 ;
     RECT  960.38 584.54 963.46 591.88 ;
     RECT  963.26 1463.6 963.74 1464.22 ;
     RECT  955.58 1312.82 964.22 1399.96 ;
     RECT  956.26 1124.24 965.18 1198.78 ;
     RECT  964.22 1312.82 965.38 1407.52 ;
     RECT  958.66 1214.12 966.14 1227.34 ;
     RECT  962.3 1240.58 966.14 1260.52 ;
     RECT  963.74 1463.6 966.14 1473.46 ;
     RECT  961.54 1094 966.34 1113.1 ;
     RECT  928.81 1574.06 966.62 1580.98 ;
     RECT  966.14 1458.98 967.58 1473.46 ;
     RECT  966.14 1214.12 967.78 1260.52 ;
     RECT  960.58 1485.86 967.78 1490.26 ;
     RECT  966.34 1105.34 968.06 1113.1 ;
     RECT  965.18 1121.72 968.06 1198.78 ;
     RECT  960.86 1272.5 968.54 1302.52 ;
     RECT  965.38 1312.82 968.54 1313.02 ;
     RECT  967.78 1214.12 969.5 1229.02 ;
     RECT  967.78 1485.86 969.5 1486.9 ;
     RECT  957.02 1501.82 970.46 1509.16 ;
     RECT  966.34 1094 970.66 1094.2 ;
     RECT  963.46 584.54 970.94 587.68 ;
     RECT  968.06 1105.34 971.14 1198.78 ;
     RECT  967.78 1240.58 971.42 1260.52 ;
     RECT  968.54 1272.5 971.42 1313.02 ;
     RECT  971.14 1132.22 971.9 1198.78 ;
     RECT  969.5 1207.4 971.9 1229.02 ;
     RECT  970.46 1501.4 972.38 1509.16 ;
     RECT  967.58 1455.2 973.06 1473.46 ;
     RECT  973.06 1456.04 973.34 1473.46 ;
     RECT  971.9 1132.22 973.54 1229.02 ;
     RECT  972.38 1501.4 973.54 1516.3 ;
     RECT  958.94 602.6 974.78 1084.54 ;
     RECT  971.9 1561.46 974.78 1561.66 ;
     RECT  959.14 1416.98 975.74 1440.7 ;
     RECT  974.78 1561.46 975.74 1562.08 ;
     RECT  975.74 1557.68 976.22 1562.08 ;
     RECT  966.62 1573.22 976.22 1580.98 ;
     RECT  975.74 1416.98 976.42 1441.54 ;
     RECT  965.38 1324.16 976.7 1407.52 ;
     RECT  973.34 1456.04 976.7 1475.14 ;
     RECT  973.54 1501.82 976.9 1516.3 ;
     RECT  971.14 1105.34 977.38 1123.18 ;
     RECT  977.38 1105.34 977.86 1121.92 ;
     RECT  976.22 1557.68 978.34 1580.98 ;
     RECT  978.34 1557.68 978.62 1562.08 ;
     RECT  977.86 1105.34 978.82 1121.5 ;
     RECT  973.54 1132.22 978.82 1228.6 ;
     RECT  922.46 -70 979 183.64 ;
     RECT  924.86 1616.06 979 1870 ;
     RECT  978.82 1105.34 979.1 1113.1 ;
     RECT  969.5 1485.44 979.78 1486.9 ;
     RECT  928.81 383.36 980.26 388.18 ;
     RECT  978.62 1557.26 980.26 1562.08 ;
     RECT  970.94 583.7 981.02 587.68 ;
     RECT  971.42 1240.58 981.02 1313.02 ;
     RECT  976.7 1322.06 981.02 1407.52 ;
     RECT  978.82 1136.84 981.7 1228.6 ;
     RECT  976.7 1456.04 982.94 1475.56 ;
     RECT  978.34 1573.22 982.94 1580.98 ;
     RECT  979.1 1103.66 983.9 1113.1 ;
     RECT  976.9 1501.82 985.34 1512.52 ;
     RECT  982.94 1453.52 986.02 1475.98 ;
     RECT  982.94 1573.22 986.02 1582.24 ;
     RECT  974.78 602.6 986.3 1090.84 ;
     RECT  983.9 1101.98 986.3 1113.1 ;
     RECT  981.7 1204.04 986.78 1228.6 ;
     RECT  981.02 1240.58 986.78 1407.52 ;
     RECT  928.81 216.2 991.19 224.8 ;
     RECT  928.81 255.26 991.19 270.16 ;
     RECT  928.81 284.24 991.19 284.44 ;
     RECT  928.81 327.5 991.19 370.96 ;
     RECT  980.26 383.36 991.19 383.98 ;
     RECT  944.26 406.46 991.19 573.82 ;
     RECT  981.02 583.7 991.19 591.88 ;
     RECT  986.3 602.6 991.19 1113.1 ;
     RECT  981.7 1136.84 991.19 1192.9 ;
     RECT  986.78 1204.04 991.19 1407.52 ;
     RECT  986.02 1453.52 991.3 1453.72 ;
     RECT  976.42 1418.24 992.06 1441.54 ;
     RECT  980.26 1557.26 992.26 1558.3 ;
     RECT  981.5 1523.66 993.02 1523.86 ;
     RECT  986.3 1535.42 993.02 1535.62 ;
     RECT  985.34 1498.46 995.62 1512.52 ;
     RECT  991.19 216.2 996.81 1407.52 ;
     RECT  979 0 997 183.64 ;
     RECT  979 1616.06 997 1800 ;
     RECT  986.02 1463.18 997.34 1475.98 ;
     RECT  979.78 1485.44 997.34 1486.06 ;
     RECT  996.81 602.6 997.54 1128.64 ;
     RECT  996.81 584.12 998.02 591.88 ;
     RECT  993.02 1523.66 998.02 1535.62 ;
     RECT  986.02 1574.06 998.3 1582.24 ;
     RECT  997.54 602.6 998.5 622.96 ;
     RECT  997.54 632.42 998.5 1128.64 ;
     RECT  996.81 1209.5 998.5 1407.52 ;
     RECT  998.02 1535.42 998.5 1535.62 ;
     RECT  998.5 632.42 998.98 1124.44 ;
     RECT  995.62 1498.46 998.98 1505.38 ;
     RECT  998.5 1211.18 999.26 1407.52 ;
     RECT  992.06 1417.82 999.26 1441.54 ;
     RECT  998.02 584.12 999.94 584.74 ;
     RECT  996.81 1137.26 999.94 1161.82 ;
     RECT  997.34 1463.18 1000.7 1486.06 ;
     RECT  998.98 1025.12 1001.38 1124.44 ;
     RECT  999.26 1211.18 1001.38 1441.54 ;
     RECT  998.98 1498.46 1001.86 1504.96 ;
     RECT  992.26 1558.1 1001.86 1558.3 ;
     RECT  998.3 1569.44 1003.58 1582.24 ;
     RECT  996.81 406.46 1003.78 573.82 ;
     RECT  1003.58 1565.24 1003.78 1582.24 ;
     RECT  1003.78 406.46 1004.52 561.22 ;
     RECT  998.98 632.42 1004.52 1016.08 ;
     RECT  1001.38 1212.86 1004.54 1441.54 ;
     RECT  1004.52 794.44 1004.74 1016.08 ;
     RECT  999.94 1147.76 1004.74 1161.82 ;
     RECT  1004.52 726.04 1005.22 757.78 ;
     RECT  998.02 1523.66 1005.7 1523.86 ;
     RECT  1000.7 1460.24 1005.98 1486.06 ;
     RECT  1004.52 632.42 1006.18 713.26 ;
     RECT  1005.22 755.48 1006.66 757.78 ;
     RECT  996.81 1171.28 1006.66 1200.88 ;
     RECT  1001.38 1080.56 1007.14 1124.44 ;
     RECT  1003.78 571.52 1007.42 573.82 ;
     RECT  1007.42 571.52 1007.62 574.66 ;
     RECT  1004.54 1212.86 1007.62 1445.32 ;
     RECT  1005.98 1460.24 1007.62 1488.16 ;
     RECT  1001.38 1025.12 1008.1 1071.94 ;
     RECT  1007.14 1080.56 1008.1 1121.08 ;
     RECT  1006.66 1171.28 1008.1 1192.9 ;
     RECT  1007.62 1339.7 1008.1 1441.54 ;
     RECT  1007.62 573.2 1008.58 574.66 ;
     RECT  1004.52 445.6 1008.785 462.48 ;
     RECT  1004.52 514 1008.785 530.88 ;
     RECT  1005.22 726.04 1008.785 745.18 ;
     RECT  1004.74 794.44 1008.785 1000.12 ;
     RECT  999.94 584.54 1008.86 584.74 ;
     RECT  1004.52 406.46 1008.92 426.75 ;
     RECT  1004.52 546.73 1008.92 561.22 ;
     RECT  1006.18 632.42 1008.92 708.65 ;
     RECT  1007.62 1212.86 1009.06 1328.98 ;
     RECT  1008.1 1395.56 1009.06 1441.54 ;
     RECT  1004.74 1011.68 1009.34 1016.08 ;
     RECT  1008.1 1025.12 1009.34 1071.52 ;
     RECT  1003.78 1565.24 1009.54 1565.44 ;
     RECT  1004.74 1154.9 1009.82 1161.82 ;
     RECT  1008.785 794.44 1010.02 800.62 ;
     RECT  1007.62 1463.6 1010.5 1488.16 ;
     RECT  998.5 602.6 1010.78 602.8 ;
     RECT  998.5 615.62 1010.78 622.96 ;
     RECT  1010.5 1485.44 1010.78 1488.16 ;
     RECT  1001.86 1498.46 1010.78 1504.54 ;
     RECT  1008.785 445.6 1011.385 451.08 ;
     RECT  1008.785 514 1011.385 527.62 ;
     RECT  1008.785 726.04 1011.385 731.52 ;
     RECT  1010.02 794.44 1011.385 799.92 ;
     RECT  1008.92 406.46 1011.52 424.15 ;
     RECT  1008.92 632.42 1011.52 706.05 ;
     RECT  1003.78 1574.06 1011.94 1582.24 ;
     RECT  997 -70 1012.7 183.64 ;
     RECT  1011.94 1574.06 1012.9 1577.2 ;
     RECT  1008.86 584.54 1013.18 586.84 ;
     RECT  1006.66 756.74 1013.18 757.78 ;
     RECT  1008.785 810.5 1013.18 1000.12 ;
     RECT  1009.34 1011.68 1013.18 1071.52 ;
     RECT  1013.18 584.54 1013.66 588.94 ;
     RECT  1010.78 602.6 1013.66 622.96 ;
     RECT  1008.92 546.74 1013.86 561.22 ;
     RECT  1008.785 743.3 1014.14 745.18 ;
     RECT  1009.82 1154.9 1014.34 1162.66 ;
     RECT  1009.06 1212.86 1014.62 1272.7 ;
     RECT  1011.385 524.9 1014.82 527.62 ;
     RECT  1013.86 556.4 1015.1 561.22 ;
     RECT  1014.14 743.3 1015.1 748.12 ;
     RECT  1013.18 756.74 1015.1 763.24 ;
     RECT  1008.1 1171.7 1015.1 1192.9 ;
     RECT  1010.78 1485.44 1015.1 1504.54 ;
     RECT  1011.52 632.42 1015.3 702.76 ;
     RECT  1013.18 810.5 1015.3 1071.52 ;
     RECT  1015.1 1171.7 1015.58 1193.32 ;
     RECT  1015.3 810.5 1016.26 810.7 ;
     RECT  1009.06 1395.56 1016.74 1440.28 ;
     RECT  1015.1 1485.44 1016.74 1512.94 ;
     RECT  1015.1 575.72 1017.02 575.92 ;
     RECT  1013.66 584.54 1017.02 622.96 ;
     RECT  1008.1 1085.6 1017.02 1121.08 ;
     RECT  1009.06 1282.16 1017.5 1328.98 ;
     RECT  1008.1 1339.7 1017.5 1386.52 ;
     RECT  1012.7 1454.78 1017.5 1454.98 ;
     RECT  1010.5 1463.6 1017.5 1474.3 ;
     RECT  1012.9 1574.06 1017.5 1574.26 ;
     RECT  1011.385 796.64 1017.7 799.36 ;
     RECT  1017.5 1282.16 1017.7 1386.52 ;
     RECT  1014.82 527.42 1017.98 527.62 ;
     RECT  1017.7 1312.82 1018.46 1386.52 ;
     RECT  1016.74 1395.56 1018.46 1438.18 ;
     RECT  1015.3 822.26 1018.94 1071.52 ;
     RECT  1015.1 743.3 1019.9 763.24 ;
     RECT  1004.52 775.64 1019.9 785.08 ;
     RECT  1017.98 527.42 1020.58 534.76 ;
     RECT  1015.58 1171.7 1020.86 1196.26 ;
     RECT  1014.62 1206.98 1020.86 1272.7 ;
     RECT  1013.86 546.74 1021.34 546.94 ;
     RECT  1017.5 1454.78 1021.34 1474.3 ;
     RECT  1016.74 1485.44 1021.34 1490.68 ;
     RECT  996.81 383.78 1021.54 383.98 ;
     RECT  1019.9 743.3 1022.3 785.08 ;
     RECT  1017.02 1085.6 1022.3 1124.44 ;
     RECT  999.94 1137.26 1022.3 1137.46 ;
     RECT  1014.34 1161.62 1022.3 1162.66 ;
     RECT  1020.86 1171.7 1022.3 1272.7 ;
     RECT  1017.7 1282.16 1022.3 1303.36 ;
     RECT  1022.3 1161.62 1022.5 1272.7 ;
     RECT  1022.3 1085.6 1022.78 1140.4 ;
     RECT  1018.94 822.26 1023.26 1074.46 ;
     RECT  1022.78 1083.08 1023.26 1140.4 ;
     RECT  1021.34 538.76 1023.46 546.94 ;
     RECT  1016.06 1524.5 1023.74 1524.7 ;
     RECT  1020.58 527.42 1023.94 527.62 ;
     RECT  1023.46 538.76 1024.42 538.96 ;
     RECT  1018.46 1312.82 1024.42 1438.18 ;
     RECT  1017.7 796.64 1024.7 796.84 ;
     RECT  1023.26 822.26 1024.9 1140.4 ;
     RECT  1024.42 1410.26 1025.18 1438.18 ;
     RECT  996.81 216.2 1025.86 224.8 ;
     RECT  1022.3 736.16 1025.86 785.08 ;
     RECT  1024.9 822.26 1026.34 1137.46 ;
     RECT  1017.5 1565.66 1026.34 1574.26 ;
     RECT  1024.7 795.8 1026.62 796.84 ;
     RECT  1026.34 822.26 1026.82 1074.88 ;
     RECT  1026.34 1569.02 1027.78 1569.64 ;
     RECT  1016.74 1499.3 1028.06 1512.94 ;
     RECT  1026.62 795.8 1028.26 803.14 ;
     RECT  1025.86 739.1 1028.74 785.08 ;
     RECT  1026.34 1089.38 1028.74 1137.46 ;
     RECT  1022.5 1161.62 1028.74 1272.28 ;
     RECT  1017.02 575.72 1029.5 622.96 ;
     RECT  1015.3 640.82 1029.7 702.76 ;
     RECT  1026.82 822.26 1029.98 1071.94 ;
     RECT  996.81 284.24 1030.66 284.44 ;
     RECT  1028.74 1211.6 1030.66 1272.28 ;
     RECT  1029.5 571.94 1030.94 622.96 ;
     RECT  1028.74 739.1 1031.62 784.24 ;
     RECT  1031.62 739.1 1032.1 760.3 ;
     RECT  1021.82 1151.54 1032.1 1151.74 ;
     RECT  1027.78 1569.44 1032.1 1569.64 ;
     RECT  1031.62 769.76 1032.58 784.24 ;
     RECT  1023.74 1524.5 1032.58 1527.64 ;
     RECT  1025.86 216.2 1033.06 221.86 ;
     RECT  1032.58 1524.5 1033.54 1524.7 ;
     RECT  1015.1 556.4 1033.82 561.64 ;
     RECT  1033.06 216.2 1034.02 221.44 ;
     RECT  1028.74 1101.98 1034.02 1137.46 ;
     RECT  1028.26 802.94 1034.5 803.14 ;
     RECT  1034.02 1124.24 1034.5 1137.46 ;
     RECT  996.81 327.5 1034.98 370.96 ;
     RECT  1032.58 769.76 1035.46 783.4 ;
     RECT  1034.02 1101.98 1035.46 1113.1 ;
     RECT  1029.98 815.12 1035.74 1071.94 ;
     RECT  1021.34 1454.78 1035.94 1490.68 ;
     RECT  1035.74 815.12 1036.22 1074.46 ;
     RECT  1024.42 1312.82 1036.42 1399.96 ;
     RECT  1032.1 739.1 1036.7 759.46 ;
     RECT  1011.52 406.46 1036.9 421.78 ;
     RECT  1033.82 553.04 1036.9 561.64 ;
     RECT  1035.46 770.18 1036.9 783.4 ;
     RECT  1028.74 1161.62 1036.9 1199.2 ;
     RECT  996.81 255.26 1037.38 270.16 ;
     RECT  1036.22 806.72 1037.86 1074.46 ;
     RECT  1036.42 1312.82 1037.86 1395.76 ;
     RECT  1036.9 1161.62 1038.62 1163.08 ;
     RECT  1030.66 1212.86 1038.62 1272.28 ;
     RECT  1022.3 1281.74 1038.62 1303.36 ;
     RECT  1036.7 737.42 1038.82 759.46 ;
     RECT  1037.86 806.72 1038.82 1073.2 ;
     RECT  1034.5 1132.22 1038.82 1137.46 ;
     RECT  1029.7 644.18 1039.3 702.76 ;
     RECT  1036.9 776.48 1039.3 783.4 ;
     RECT  1035.46 1101.98 1039.3 1102.18 ;
     RECT  1028.74 1091.48 1039.58 1091.68 ;
     RECT  1038.82 863.42 1039.78 1073.2 ;
     RECT  1030.94 571.94 1040.06 630.1 ;
     RECT  1040.06 571.94 1040.26 632.62 ;
     RECT  1025.18 1410.26 1040.26 1444.48 ;
     RECT  997 1616.06 1040.26 1870 ;
     RECT  1035.94 1458.56 1040.54 1490.68 ;
     RECT  1028.06 1499.3 1040.54 1514.2 ;
     RECT  1040.54 1458.56 1041.02 1514.2 ;
     RECT  1037.18 1524.08 1041.02 1524.28 ;
     RECT  1036.9 406.46 1041.7 421.36 ;
     RECT  1038.62 1212.86 1042.46 1303.36 ;
     RECT  1038.82 806.72 1042.94 854.8 ;
     RECT  1039.58 1091.48 1043.14 1098.82 ;
     RECT  1042.94 805.88 1044.1 854.8 ;
     RECT  1040.26 1410.26 1044.1 1441.12 ;
     RECT  1036.9 556.4 1044.58 561.64 ;
     RECT  1044.1 1410.26 1044.58 1439.44 ;
     RECT  1034.98 327.5 1045.06 349.12 ;
     RECT  1036.9 1175.9 1045.34 1199.2 ;
     RECT  1042.46 1208.66 1045.34 1303.36 ;
     RECT  1034.98 363.62 1045.54 370.96 ;
     RECT  1045.34 1175.9 1045.54 1303.36 ;
     RECT  1039.3 660.56 1046.02 702.76 ;
     RECT  1037.86 1319.54 1046.02 1395.76 ;
     RECT  1044.1 805.88 1046.3 809.02 ;
     RECT  1044.1 822.26 1046.5 854.8 ;
     RECT  1039.78 1006.22 1046.5 1073.2 ;
     RECT  1045.54 1175.9 1046.5 1208.86 ;
     RECT  1039.3 644.18 1046.98 651.94 ;
     RECT  1039.3 776.48 1046.98 780.46 ;
     RECT  1041.02 1458.56 1046.98 1524.28 ;
     RECT  1035.46 1112.06 1047.26 1113.1 ;
     RECT  1046.5 838.22 1047.46 854.8 ;
     RECT  1038.82 1137.26 1047.74 1137.46 ;
     RECT  1041.7 406.46 1047.94 407.08 ;
     RECT  1046.02 1392.62 1047.94 1395.76 ;
     RECT  1047.74 1137.26 1048.22 1143.34 ;
     RECT  1037.38 262.82 1048.42 270.16 ;
     RECT  1046.5 1006.22 1048.42 1011.88 ;
     RECT  1048.22 1130.96 1048.42 1143.34 ;
     RECT  1044.58 1410.26 1048.42 1438.6 ;
     RECT  1012.7 1603.04 1048.42 1603.24 ;
     RECT  1039.78 863.42 1048.9 997.18 ;
     RECT  1046.5 1175.9 1048.9 1198.78 ;
     RECT  1048.42 1006.22 1049.38 1006.42 ;
     RECT  1040.26 571.94 1049.86 622.96 ;
     RECT  1048.42 1130.96 1050.34 1137.46 ;
     RECT  1040.26 632.42 1050.62 632.62 ;
     RECT  1050.62 632.42 1050.82 640.6 ;
     RECT  1048.9 1175.9 1051.1 1193.32 ;
     RECT  1045.54 363.62 1051.3 363.82 ;
     RECT  1046.3 800 1051.3 809.02 ;
     RECT  1046.5 1208.24 1051.3 1208.86 ;
     RECT  1048.42 1410.26 1051.3 1412.14 ;
     RECT  1046.02 1319.54 1051.58 1382.32 ;
     RECT  1038.82 738.68 1051.78 759.46 ;
     RECT  1046.98 777.32 1052.54 780.46 ;
     RECT  1041.7 416.54 1053.22 421.36 ;
     RECT  1046.5 1025.12 1053.22 1073.2 ;
     RECT  1051.58 1317.86 1053.7 1382.32 ;
     RECT  1047.26 1081.82 1053.98 1082.02 ;
     RECT  1051.3 800 1054.18 800.2 ;
     RECT  1047.26 1112.06 1054.46 1116.46 ;
     RECT  1044.58 556.4 1054.66 561.22 ;
     RECT  1051.3 1410.26 1054.66 1411.72 ;
     RECT  1051.3 808.82 1054.94 809.02 ;
     RECT  1046.5 822.26 1054.94 828.76 ;
     RECT  1046.98 1458.56 1055.42 1474.3 ;
     RECT  1046.98 1485.02 1055.42 1524.28 ;
     RECT  1049.86 583.28 1055.62 622.96 ;
     RECT  1050.62 1101.98 1055.62 1102.18 ;
     RECT  1055.42 1458.56 1055.62 1524.28 ;
     RECT  1046.02 662.66 1056.1 702.76 ;
     RECT  1053.22 416.54 1056.58 420.1 ;
     RECT  1055.62 1497.2 1057.34 1524.28 ;
     RECT  1051.78 742.88 1058.02 759.46 ;
     RECT  1053.98 1081.82 1058.02 1082.86 ;
     RECT  1049.86 571.94 1058.3 572.98 ;
     RECT  1055.62 583.28 1058.3 588.1 ;
     RECT  1055.62 598.4 1058.3 622.96 ;
     RECT  1051.3 1208.66 1058.3 1208.86 ;
     RECT  1058.3 571.94 1058.5 588.1 ;
     RECT  1058.02 743.72 1058.5 759.46 ;
     RECT  1058.02 1081.82 1058.5 1082.02 ;
     RECT  1038.62 1159.94 1058.5 1163.08 ;
     RECT  1054.94 808.82 1058.78 828.76 ;
     RECT  1047.46 841.16 1058.78 854.8 ;
     RECT  1048.42 1420.76 1058.78 1438.6 ;
     RECT  1052.54 777.32 1059.26 782.98 ;
     RECT  1058.78 808.82 1059.74 854.8 ;
     RECT  1048.9 867.62 1059.74 997.18 ;
     RECT  1059.74 808.82 1059.94 997.18 ;
     RECT  1058.5 744.14 1060.22 759.46 ;
     RECT  1054.46 1111.64 1060.22 1116.46 ;
     RECT  1058.5 1161.62 1060.22 1163.08 ;
     RECT  1051.1 1173.8 1060.22 1193.32 ;
     RECT  1058.3 1208.66 1060.22 1209.28 ;
     RECT  1045.54 1217.9 1060.22 1303.36 ;
     RECT  1058.78 1420.76 1060.42 1440.28 ;
     RECT  1059.26 775.64 1061.18 782.98 ;
     RECT  1059.94 808.82 1061.18 829.6 ;
     RECT  1060.22 1217.9 1061.18 1304.2 ;
     RECT  1053.7 1317.86 1061.18 1378.12 ;
     RECT  1056.1 664.34 1061.38 702.76 ;
     RECT  1061.18 807.14 1061.38 829.6 ;
     RECT  1015.58 1548.86 1061.38 1549.06 ;
     RECT  1060.22 1161.62 1061.86 1195.84 ;
     RECT  1061.18 775.64 1062.14 788.44 ;
     RECT  1055.62 1458.56 1062.14 1488.16 ;
     RECT  1062.14 775.64 1062.34 788.86 ;
     RECT  1061.38 807.14 1062.62 828.76 ;
     RECT  1060.22 1207.4 1062.62 1209.28 ;
     RECT  1061.18 1217.9 1062.62 1378.12 ;
     RECT  1056.58 416.54 1062.82 418 ;
     RECT  1048.42 269.96 1063.3 270.16 ;
     RECT  1062.14 1451.42 1063.3 1488.16 ;
     RECT  1057.34 1497.2 1063.3 1528.06 ;
     RECT  1060.22 744.14 1063.58 765.34 ;
     RECT  1060.22 1104.5 1063.58 1116.46 ;
     RECT  1053.22 1031.84 1063.78 1073.2 ;
     RECT  1061.38 677.78 1064.26 702.76 ;
     RECT  1063.3 1451.42 1064.74 1481.86 ;
     RECT  1062.62 1207.4 1065.22 1378.12 ;
     RECT  1063.3 1526.18 1065.5 1528.06 ;
     RECT  1062.82 416.54 1065.7 416.74 ;
     RECT  1064.26 677.78 1066.66 681.76 ;
     RECT  1060.42 1420.76 1066.94 1436.92 ;
     RECT  1012.7 -70 1067 184.06 ;
     RECT  1040.26 1622 1067 1870 ;
     RECT  1058.3 598.4 1067.42 627.16 ;
     RECT  1061.38 664.34 1067.62 664.96 ;
     RECT  1063.78 1031.84 1067.62 1071.94 ;
     RECT  1064.74 1451.42 1067.62 1478.5 ;
     RECT  1061.86 1161.62 1067.9 1181.56 ;
     RECT  1064.26 693.32 1068.1 702.76 ;
     RECT  1054.66 561.02 1068.38 561.22 ;
     RECT  1063.58 744.14 1068.86 766.6 ;
     RECT  1063.58 1104.5 1068.86 1124.86 ;
     RECT  1050.34 1137.26 1068.86 1137.46 ;
     RECT  1066.94 1420.34 1068.86 1436.92 ;
     RECT  438.14 197.72 1069.06 197.92 ;
     RECT  1063.3 1497.2 1069.34 1516.3 ;
     RECT  1045.06 341.78 1069.54 349.12 ;
     RECT  1062.62 805.46 1069.54 828.76 ;
     RECT  1067.9 1159.52 1069.54 1181.56 ;
     RECT  1068.86 1420.34 1070.02 1438.6 ;
     RECT  1069.54 806.72 1070.3 828.76 ;
     RECT  1059.94 840.74 1070.3 997.18 ;
     RECT  1054.66 1411.52 1070.3 1411.72 ;
     RECT  1070.02 1420.34 1070.3 1437.76 ;
     RECT  1050.82 640.4 1070.5 640.6 ;
     RECT  1069.34 1493.84 1070.5 1516.3 ;
     RECT  1062.34 788.24 1071.26 788.86 ;
     RECT  1069.54 1165.82 1071.26 1181.56 ;
     RECT  1061.86 1192.7 1071.26 1195.84 ;
     RECT  1067.42 598.4 1072.22 629.26 ;
     RECT  1071.74 731.12 1072.22 731.32 ;
     RECT  1071.26 788.24 1072.22 790.96 ;
     RECT  1071.26 1165.82 1072.42 1195.84 ;
     RECT  1068.38 554.72 1072.7 561.22 ;
     RECT  1072.22 788.24 1072.7 791.8 ;
     RECT  1067.62 1065.02 1072.7 1071.94 ;
     RECT  1067.62 1031.84 1072.9 1054.3 ;
     RECT  1072.42 1165.82 1072.9 1176.1 ;
     RECT  1072.42 1188.5 1072.9 1195.84 ;
     RECT  1062.34 775.64 1073.18 777.1 ;
     RECT  1072.7 788.24 1073.18 792.22 ;
     RECT  1047.94 406.46 1073.38 406.66 ;
     RECT  1065.22 1209.92 1073.38 1378.12 ;
     RECT  1068.86 743.3 1073.66 766.6 ;
     RECT  1073.18 775.64 1073.66 792.22 ;
     RECT  1068.1 695 1073.86 702.76 ;
     RECT  1072.7 1022.18 1073.86 1023.22 ;
     RECT  1043.14 1091.48 1074.14 1091.68 ;
     RECT  1072.7 554.72 1074.34 562.48 ;
     RECT  1046.98 651.74 1074.34 651.94 ;
     RECT  1058.5 572.78 1074.62 578.44 ;
     RECT  1072.9 1189.76 1074.62 1195.84 ;
     RECT  1073.38 1209.92 1074.62 1210.12 ;
     RECT  1074.62 571.94 1075.1 578.44 ;
     RECT  1058.5 587.06 1075.1 588.1 ;
     RECT  1070.5 1516.1 1075.1 1516.3 ;
     RECT  1065.5 1526.18 1075.1 1531.84 ;
     RECT  1075.1 1516.1 1075.3 1531.84 ;
     RECT  1071.26 1565.24 1075.3 1565.44 ;
     RECT  1072.22 598.4 1075.58 629.68 ;
     RECT  1068.86 1104.5 1075.58 1137.46 ;
     RECT  1074.34 561.02 1075.78 562.48 ;
     RECT  1073.66 743.3 1075.78 792.22 ;
     RECT  1070.3 1411.52 1075.78 1437.76 ;
     RECT  1073.86 695 1076.26 696.88 ;
     RECT  1075.78 1411.52 1078.18 1429.78 ;
     RECT  1075.58 1104.5 1078.94 1145.86 ;
     RECT  1072.22 1155.32 1078.94 1155.52 ;
     RECT  1070.5 1493.84 1078.94 1504.96 ;
     RECT  1075.3 1531.64 1079.14 1531.84 ;
     RECT  1070.3 806.72 1079.42 997.18 ;
     RECT  1076.06 1447.22 1079.42 1447.42 ;
     RECT  1067.62 1456.04 1079.42 1478.5 ;
     RECT  1075.58 598.4 1079.62 630.1 ;
     RECT  1072.7 1065.02 1079.9 1073.2 ;
     RECT  1076.26 696.68 1080.1 696.88 ;
     RECT  1079.62 598.4 1080.38 608.26 ;
     RECT  1078.94 1104.5 1080.38 1155.52 ;
     RECT  1075.78 775.64 1080.86 792.22 ;
     RECT  1079.42 1447.22 1081.06 1478.5 ;
     RECT  1066.66 677.78 1081.34 680.5 ;
     RECT  1072.9 1170.86 1081.34 1176.1 ;
     RECT  1078.94 1493.84 1081.54 1505.38 ;
     RECT  1075.78 561.02 1082.02 561.22 ;
     RECT  1080.86 775.64 1082.3 796 ;
     RECT  1079.42 806.72 1082.3 1004.74 ;
     RECT  1052.06 230.48 1082.5 230.68 ;
     RECT  1072.9 1032.68 1082.78 1054.3 ;
     RECT  1079.9 1065.02 1082.78 1075.72 ;
     RECT  1082.78 1032.68 1083.26 1075.72 ;
     RECT  1074.14 1086.44 1083.26 1091.68 ;
     RECT  1074.62 1189.76 1083.26 1210.12 ;
     RECT  1034.02 221.24 1083.46 221.44 ;
     RECT  1081.06 1447.22 1083.46 1473.88 ;
     RECT  1079.62 617.72 1083.74 630.1 ;
     RECT  1069.54 348.92 1083.94 349.12 ;
     RECT  1081.34 1170.86 1084.22 1177.36 ;
     RECT  1083.26 1186.4 1084.22 1210.12 ;
     RECT  1081.54 1493.84 1084.22 1504.96 ;
     RECT  1083.74 617.72 1084.42 635.56 ;
     RECT  1084.42 626.96 1084.7 635.56 ;
     RECT  1077.02 644.18 1084.7 644.38 ;
     RECT  1067 0 1085 184.06 ;
     RECT  1067 1622 1085 1800 ;
     RECT  1075.1 571.94 1085.18 588.1 ;
     RECT  1083.26 712.64 1085.38 712.84 ;
     RECT  1073.38 1218.74 1085.38 1378.12 ;
     RECT  1085.18 569.84 1085.66 588.1 ;
     RECT  1080.38 597.56 1085.66 608.26 ;
     RECT  1078.18 1411.52 1085.86 1429.36 ;
     RECT  1085.86 1414.04 1086.34 1421.8 ;
     RECT  1083.46 1447.22 1086.62 1471.78 ;
     RECT  1084.7 626.96 1086.82 644.38 ;
     RECT  1067.62 664.76 1087.3 664.96 ;
     RECT  1084.22 1170.86 1087.3 1210.12 ;
     RECT  1085.38 1263.26 1087.3 1378.12 ;
     RECT  1084.22 1483.34 1087.3 1504.96 ;
     RECT  1075.3 1516.1 1087.3 1520.08 ;
     RECT  1086.82 626.96 1087.78 635.56 ;
     RECT  1086.34 1414.04 1087.78 1420.54 ;
     RECT  1086.62 1438.82 1087.78 1471.78 ;
     RECT  1081.34 677.78 1088.26 683.86 ;
     RECT  1083.26 1032.68 1088.26 1091.68 ;
     RECT  1087.3 1172.96 1088.26 1210.12 ;
     RECT  1087.3 1270.82 1088.26 1378.12 ;
     RECT  1086.82 644.18 1088.74 644.38 ;
     RECT  1082.3 775.64 1088.74 1004.74 ;
     RECT  1087.78 1448.9 1088.74 1471.36 ;
     RECT  1087.78 629.9 1089.22 635.56 ;
     RECT  1087.78 1438.82 1089.22 1439.02 ;
     RECT  1087.3 1516.1 1089.22 1516.3 ;
     RECT  1085.66 569.84 1089.5 608.26 ;
     RECT  1084.42 617.72 1089.5 617.92 ;
     RECT  1075.78 743.3 1089.5 766.18 ;
     RECT  1088.74 775.64 1089.5 790.96 ;
     RECT  1085.38 1218.74 1089.7 1254.64 ;
     RECT  1088.26 1032.68 1090.18 1074.88 ;
     RECT  1089.7 1219.16 1090.18 1254.64 ;
     RECT  1085 -70 1090.66 184.06 ;
     RECT  1088.26 1172.96 1090.66 1206.34 ;
     RECT  1045.06 327.5 1091.14 327.7 ;
     RECT  1088.74 1448.9 1091.14 1453.3 ;
     RECT  1088.74 1463.18 1092.1 1471.36 ;
     RECT  1089.5 569.84 1093.06 617.92 ;
     RECT  1090.18 1032.68 1093.06 1060.18 ;
     RECT  1088.26 1083.92 1093.06 1091.68 ;
     RECT  1087.3 1489.22 1093.06 1504.96 ;
     RECT  1088.74 799.58 1094.5 1004.74 ;
     RECT  1093.06 1032.68 1094.5 1058.5 ;
     RECT  1091.14 1448.9 1095.46 1449.1 ;
     RECT  1089.5 743.3 1095.94 790.96 ;
     RECT  1095.74 1018.82 1096.42 1019.02 ;
     RECT  1087.78 1420.34 1096.42 1420.54 ;
     RECT  1093.06 1495.94 1096.42 1504.96 ;
     RECT  1090.18 1074.68 1096.9 1074.88 ;
     RECT  1072.22 725.66 1097.18 731.32 ;
     RECT  1095.94 743.3 1097.18 783.4 ;
     RECT  1094.5 1032.68 1097.38 1053.04 ;
     RECT  1092.1 1468.64 1097.66 1471.36 ;
     RECT  1090.66 1172.96 1097.86 1176.1 ;
     RECT  1097.38 1032.68 1098.34 1049.68 ;
     RECT  1080.38 1104.5 1098.34 1159.72 ;
     RECT  1094.5 799.58 1099.3 997.18 ;
     RECT  1088.26 1270.82 1099.3 1377.7 ;
     RECT  1090.66 1186.4 1099.78 1206.34 ;
     RECT  1099.3 1270.82 1100.26 1279.84 ;
     RECT  1093.06 569.84 1100.54 610.78 ;
     RECT  1090.18 1219.16 1101.02 1252.96 ;
     RECT  1099.78 1187.66 1101.22 1206.34 ;
     RECT  1100.26 1271.24 1101.22 1279.84 ;
     RECT  1100.54 565.22 1101.5 610.78 ;
     RECT  1098.34 1032.68 1101.7 1038.34 ;
     RECT  1101.22 1187.66 1101.7 1196.26 ;
     RECT  1099.3 799.58 1102.18 950.14 ;
     RECT  1097.66 1468.64 1102.66 1482.7 ;
     RECT  1088.26 677.78 1103.14 680.5 ;
     RECT  1097.18 725.66 1103.14 783.4 ;
     RECT  1102.66 1468.64 1104.58 1468.84 ;
     RECT  1101.02 1217.06 1105.06 1252.96 ;
     RECT  1097.18 1023.44 1105.82 1023.64 ;
     RECT  1101.22 1204.88 1105.82 1206.34 ;
     RECT  1096.42 1500.98 1106.02 1504.96 ;
     RECT  1089.22 635.36 1106.5 635.56 ;
     RECT  1099.3 1290.56 1106.5 1377.7 ;
     RECT  1047.94 1392.62 1106.98 1392.82 ;
     RECT  1106.02 1504.76 1106.98 1504.96 ;
     RECT  1102.18 881.48 1107.74 950.14 ;
     RECT  1099.3 958.76 1107.74 997.18 ;
     RECT  1106.5 1290.56 1107.94 1371.82 ;
     RECT  1107.74 881.48 1108.22 997.18 ;
     RECT  1107.94 1361.96 1108.42 1371.82 ;
     RECT  1077.5 546.32 1108.7 546.52 ;
     RECT  1098.34 1049.48 1108.7 1049.68 ;
     RECT  1105.82 1204.88 1108.7 1207.6 ;
     RECT  1105.06 1217.06 1108.7 1252.54 ;
     RECT  1101.22 1276.7 1108.7 1279.84 ;
     RECT  1108.7 1204.88 1108.9 1252.54 ;
     RECT  1108.42 1361.96 1108.9 1368.46 ;
     RECT  1108.9 1204.88 1109.38 1209.28 ;
     RECT  1101.5 561.86 1109.66 616.66 ;
     RECT  1108.7 540.44 1110.14 546.52 ;
     RECT  1108.9 1367.84 1110.34 1368.46 ;
     RECT  1105.82 1022.6 1111.1 1023.64 ;
     RECT  1101.7 1038.14 1111.1 1038.34 ;
     RECT  1110.34 1368.26 1111.3 1368.46 ;
     RECT  1102.18 799.58 1111.58 868.66 ;
     RECT  1108.22 881.48 1111.58 1002.22 ;
     RECT  1101.7 1187.66 1111.78 1192.9 ;
     RECT  1110.14 538.76 1112.06 546.52 ;
     RECT  1111.1 1022.6 1112.06 1038.34 ;
     RECT  1098.34 1104.5 1112.06 1155.52 ;
     RECT  1097.86 1173.8 1112.06 1176.1 ;
     RECT  1103.14 725.66 1112.54 754.84 ;
     RECT  1111.58 799.58 1112.54 1002.22 ;
     RECT  1112.06 1022.18 1112.74 1038.34 ;
     RECT  1112.54 796.64 1113.22 1002.22 ;
     RECT  1112.06 1104.5 1113.5 1162.24 ;
     RECT  1112.06 1173.8 1113.5 1177.36 ;
     RECT  1103.14 765.98 1113.98 783.4 ;
     RECT  1113.98 765.56 1115.42 783.4 ;
     RECT  1108.7 1276.7 1115.42 1281.94 ;
     RECT  1107.94 1290.56 1115.42 1347.88 ;
     RECT  1112.74 1022.18 1115.62 1026.16 ;
     RECT  1108.9 1219.16 1115.9 1252.54 ;
     RECT  1113.5 1262 1115.9 1262.2 ;
     RECT  1115.42 1276.7 1115.9 1347.88 ;
     RECT  1109.66 561.02 1116.38 616.66 ;
     RECT  1112.06 1011.68 1116.58 1011.88 ;
     RECT  1112.54 721.04 1116.86 754.84 ;
     RECT  1115.42 765.56 1116.86 783.82 ;
     RECT  1115.9 1273.34 1116.86 1347.88 ;
     RECT  1113.22 799.58 1117.34 1002.22 ;
     RECT  1116.86 1273.34 1117.34 1351.66 ;
     RECT  1112.06 534.98 1117.82 546.52 ;
     RECT  1111.78 1190.18 1117.82 1192.9 ;
     RECT  1109.38 1204.88 1117.82 1207.6 ;
     RECT  1103.14 680.3 1118.5 680.5 ;
     RECT  1116.86 721.04 1120.22 783.82 ;
     RECT  1117.82 534.14 1120.7 546.52 ;
     RECT  1117.82 1190.18 1120.7 1207.6 ;
     RECT  1108.7 1049.48 1121.18 1052.2 ;
     RECT  1117.34 1272.92 1121.18 1351.66 ;
     RECT  1120.22 721.04 1122.14 785.08 ;
     RECT  1117.34 799.58 1122.62 1004.74 ;
     RECT  1121.18 1272.5 1122.62 1351.66 ;
     RECT  1118.78 1362.38 1122.62 1362.58 ;
     RECT  1120.7 532.04 1123.1 546.52 ;
     RECT  1116.38 557.24 1123.1 616.66 ;
     RECT  1123.1 531.2 1123.58 616.66 ;
     RECT  1122.62 1272.5 1123.58 1362.58 ;
     RECT  1108.7 708.44 1124.06 708.64 ;
     RECT  1115.9 1219.16 1124.06 1262.2 ;
     RECT  1123.58 1272.5 1124.06 1363 ;
     RECT  1122.14 721.04 1124.54 788.86 ;
     RECT  1113.5 1104.5 1124.54 1177.36 ;
     RECT  1121.18 1048.64 1125.02 1052.2 ;
     RECT  1093.06 1091.48 1125.02 1091.68 ;
     RECT  1119.74 697.1 1125.98 697.3 ;
     RECT  1124.06 706.76 1125.98 708.64 ;
     RECT  1115.62 1022.6 1125.98 1026.16 ;
     RECT  1120.7 1187.66 1125.98 1207.6 ;
     RECT  1124.06 1219.16 1125.98 1363 ;
     RECT  1124.54 719.36 1126.46 788.86 ;
     RECT  1122.62 798.74 1126.46 1004.74 ;
     RECT  1125.02 1048.64 1126.46 1053.04 ;
     RECT  1125.02 1089.8 1126.46 1091.68 ;
     RECT  1124.54 1104.5 1126.46 1178.2 ;
     RECT  1123.58 531.2 1126.94 622.54 ;
     RECT  1126.46 719.36 1126.94 1004.74 ;
     RECT  1126.46 1048.22 1126.94 1053.04 ;
     RECT  1126.46 1089.8 1126.94 1178.2 ;
     RECT  1125.98 1187.66 1126.94 1363 ;
     RECT  1126.94 527.42 1127.19 622.54 ;
     RECT  1123.58 637.04 1127.19 637.24 ;
     RECT  1102.46 647.96 1127.19 648.16 ;
     RECT  1119.26 658.46 1127.19 658.66 ;
     RECT  1122.62 678.62 1127.19 678.82 ;
     RECT  1125.98 697.1 1127.19 708.64 ;
     RECT  1126.94 719.36 1127.19 1007.26 ;
     RECT  1125.98 1017.56 1127.19 1026.16 ;
     RECT  1112.74 1036.88 1127.19 1038.34 ;
     RECT  1126.94 1047.8 1127.19 1053.04 ;
     RECT  1126.94 1089.8 1127.19 1363 ;
     RECT  1127.19 215.36 1132.81 1583.92 ;
     RECT  1132.81 1298.54 1132.9 1322.26 ;
     RECT  1132.81 1332.14 1132.9 1363 ;
     RECT  1132.81 647.96 1133.38 658.66 ;
     RECT  1132.81 678.62 1133.38 678.82 ;
     RECT  1132.81 1089.8 1133.38 1262.2 ;
     RECT  1132.81 719.78 1133.86 868.66 ;
     RECT  1132.9 1332.98 1133.86 1363 ;
     RECT  1132.9 1298.54 1134.34 1320.16 ;
     RECT  1132.81 519.44 1134.82 587.68 ;
     RECT  1132.81 637.04 1134.82 637.24 ;
     RECT  1132.81 881.48 1135.3 1008.94 ;
     RECT  1133.38 1233.44 1135.3 1262.2 ;
     RECT  1135.3 1253.18 1135.78 1262.2 ;
     RECT  1134.82 553.88 1136.26 587.68 ;
     RECT  1133.86 737.84 1136.74 868.24 ;
     RECT  1132.81 1021.34 1136.74 1053.04 ;
     RECT  1135.78 1254.02 1136.74 1262.2 ;
     RECT  1133.86 1332.98 1136.74 1333.18 ;
     RECT  1132.81 605.96 1139.14 625.48 ;
     RECT  1133.86 1343.9 1140.1 1363 ;
     RECT  1136.74 755.48 1140.58 788.86 ;
     RECT  1139.14 608.06 1141.06 616.66 ;
     RECT  1134.34 1298.54 1141.54 1317.64 ;
     RECT  1133.38 1089.8 1142.5 1219.36 ;
     RECT  1142.5 1091.06 1142.78 1219.36 ;
     RECT  1141.06 608.06 1143.94 614.14 ;
     RECT  1136.74 1022.6 1143.94 1053.04 ;
     RECT  1142.78 1091.06 1144.42 1223.14 ;
     RECT  1141.54 1309.46 1144.42 1317.22 ;
     RECT  1133.86 719.78 1144.7 728.38 ;
     RECT  1136.74 737.84 1144.7 746.02 ;
     RECT  1140.58 757.16 1145.18 788.86 ;
     RECT  1136.74 797.9 1145.18 868.24 ;
     RECT  1145.18 757.16 1145.66 868.24 ;
     RECT  1144.42 1164.56 1145.86 1223.14 ;
     RECT  1143.94 1022.6 1146.14 1052.2 ;
     RECT  1132.81 1078.88 1146.34 1079.08 ;
     RECT  1132.81 697.1 1146.62 697.3 ;
     RECT  1135.3 980.6 1146.62 1008.94 ;
     RECT  1146.14 1021.34 1146.62 1052.2 ;
     RECT  1143.94 613.94 1146.82 614.14 ;
     RECT  1139.14 625.28 1146.82 625.48 ;
     RECT  1132.81 1067.96 1147.1 1068.16 ;
     RECT  1134.82 519.44 1147.3 542.74 ;
     RECT  1146.62 980.6 1147.3 1052.2 ;
     RECT  1135.3 881.48 1147.58 969.88 ;
     RECT  1147.3 980.6 1147.58 1008.94 ;
     RECT  1144.7 719.78 1148.54 746.02 ;
     RECT  1145.66 757.16 1149.22 871.6 ;
     RECT  1147.3 1021.34 1149.7 1050.1 ;
     RECT  1136.26 558.92 1150.66 587.68 ;
     RECT  1133.38 652.16 1151.14 658.66 ;
     RECT  1141.54 1298.54 1151.42 1300.42 ;
     RECT  1144.42 1309.46 1151.42 1310.08 ;
     RECT  1145.86 1164.56 1151.62 1200.04 ;
     RECT  1145.86 1210.76 1151.62 1223.14 ;
     RECT  1147.58 881.48 1152.1 1008.94 ;
     RECT  1136.74 1260.32 1152.1 1262.2 ;
     RECT  1132.81 1272.5 1152.38 1279 ;
     RECT  1146.62 697.1 1152.58 704.86 ;
     RECT  1151.42 1298.54 1152.58 1310.08 ;
     RECT  1152.38 1329.2 1152.86 1329.4 ;
     RECT  1151.62 1164.56 1153.06 1199.62 ;
     RECT  1152.1 1262 1153.34 1262.2 ;
     RECT  1152.38 1272.5 1153.34 1286.98 ;
     RECT  1152.58 697.1 1153.54 697.3 ;
     RECT  1135.3 1233.44 1153.54 1242.04 ;
     RECT  1152.58 1298.54 1153.54 1306.72 ;
     RECT  1140.1 1346 1153.54 1363 ;
     RECT  1148.54 719.78 1154.3 747.7 ;
     RECT  1149.22 757.16 1154.3 867.82 ;
     RECT  1153.34 1262 1154.98 1286.98 ;
     RECT  1090.66 -70 1155 178 ;
     RECT  1085 1622 1155 1870 ;
     RECT  1153.54 1346 1155.26 1360.48 ;
     RECT  1153.06 1171.28 1155.46 1199.62 ;
     RECT  1155.26 1344.32 1155.46 1360.48 ;
     RECT  1147.3 519.44 1155.74 542.32 ;
     RECT  1154.3 719.78 1155.94 867.82 ;
     RECT  1144.42 1091.06 1156.22 1155.1 ;
     RECT  1155.94 720.2 1156.42 867.82 ;
     RECT  1156.22 1090.64 1156.42 1155.1 ;
     RECT  1152.1 885.26 1156.7 1008.94 ;
     RECT  1149.7 1021.34 1156.7 1026.58 ;
     RECT  1152.86 1325 1156.7 1329.4 ;
     RECT  1155.46 1190.18 1157.38 1199.62 ;
     RECT  1153.54 1234.28 1157.38 1242.04 ;
     RECT  1155.46 1355.66 1158.34 1360.48 ;
     RECT  1156.7 1317.44 1158.82 1329.4 ;
     RECT  1155.46 1344.32 1158.82 1346.2 ;
     RECT  1158.34 1356.08 1158.82 1360.48 ;
     RECT  1155.74 519.44 1159.1 549.46 ;
     RECT  1150.66 558.92 1159.1 559.12 ;
     RECT  1150.66 569.84 1159.1 587.68 ;
     RECT  1149.7 1037.3 1159.1 1050.1 ;
     RECT  1149.02 1079.3 1159.1 1079.5 ;
     RECT  1154.98 1271.66 1159.1 1286.98 ;
     RECT  1153.54 1298.54 1159.1 1300.42 ;
     RECT  1159.1 1079.3 1159.3 1080.76 ;
     RECT  1155.46 1171.28 1159.3 1177.36 ;
     RECT  1151.62 1210.76 1159.3 1219.36 ;
     RECT  1154.98 1262 1159.3 1262.2 ;
     RECT  1158.82 1317.44 1159.3 1328.98 ;
     RECT  1159.1 1271.66 1159.78 1300.42 ;
     RECT  1159.3 1320.8 1159.78 1328.98 ;
     RECT  1156.7 885.26 1160.06 1026.58 ;
     RECT  1159.1 1037.3 1160.06 1058.5 ;
     RECT  1156.42 720.2 1160.74 746.02 ;
     RECT  1158.82 1356.08 1160.74 1359.22 ;
     RECT  1159.1 519.44 1161.98 559.12 ;
     RECT  1159.1 569.84 1161.98 591.04 ;
     RECT  1157.38 1241.84 1162.46 1242.04 ;
     RECT  1159.1 1251.08 1162.46 1251.28 ;
     RECT  1156.42 757.16 1163.42 867.82 ;
     RECT  1163.42 757.16 1163.62 871.6 ;
     RECT  1160.06 885.26 1164.38 1058.5 ;
     RECT  1147.1 1067.96 1164.38 1069.42 ;
     RECT  1163.62 827.3 1165.06 871.6 ;
     RECT  1161.98 708.44 1165.54 708.64 ;
     RECT  1162.46 1241.84 1166.3 1251.28 ;
     RECT  1159.78 1320.8 1166.5 1322.68 ;
     RECT  1160.74 727.76 1167.26 746.02 ;
     RECT  1163.62 757.16 1167.26 818.68 ;
     RECT  1158.82 1346 1167.26 1346.2 ;
     RECT  1159.78 1286.36 1167.46 1300.42 ;
     RECT  1159.3 1174.22 1168.22 1177.36 ;
     RECT  1164.38 885.26 1168.7 1069.42 ;
     RECT  1166.3 1238.06 1168.7 1251.28 ;
     RECT  1168.7 881.48 1168.9 1069.42 ;
     RECT  1159.1 618.14 1169.18 618.34 ;
     RECT  1159.3 1219.16 1169.18 1219.36 ;
     RECT  1157.38 1192.7 1169.66 1199.62 ;
     RECT  1162.46 1310.72 1170.14 1310.92 ;
     RECT  1169.18 610.16 1170.82 618.34 ;
     RECT  1169.66 1192.7 1171.1 1200.46 ;
     RECT  1163.9 1210.34 1171.1 1210.54 ;
     RECT  1168.7 1234.7 1171.1 1252.54 ;
     RECT  1171.1 1234.7 1172.06 1252.96 ;
     RECT  1155 0 1173 178 ;
     RECT  1155 1622 1173 1800 ;
     RECT  1168.22 1170.44 1173.02 1177.36 ;
     RECT  1171.1 1192.7 1173.02 1210.54 ;
     RECT  1172.06 1234.28 1173.02 1252.96 ;
     RECT  1167.26 727.76 1173.5 818.68 ;
     RECT  1165.06 827.3 1173.5 867.82 ;
     RECT  1168.9 881.48 1173.5 977.44 ;
     RECT  1167.26 1343.48 1173.5 1346.2 ;
     RECT  1173.5 727.76 1174.66 977.44 ;
     RECT  1167.46 1286.36 1175.14 1300 ;
     RECT  1173.5 703.82 1175.62 704.02 ;
     RECT  1168.7 716.42 1175.62 716.62 ;
     RECT  1161.98 519.44 1176.1 591.04 ;
     RECT  1173.02 1233.44 1176.1 1252.96 ;
     RECT  1171.58 1325 1176.38 1325.2 ;
     RECT  1168.9 989.84 1176.86 1069.42 ;
     RECT  1174.66 934.4 1178.3 977.44 ;
     RECT  1156.42 1090.64 1178.5 1153.42 ;
     RECT  1176.1 519.86 1179.74 591.04 ;
     RECT  1174.66 727.76 1179.94 924.94 ;
     RECT  1176.86 989.84 1180.42 1069.84 ;
     RECT  1176.38 1325 1180.7 1332.34 ;
     RECT  1173.5 1343.48 1180.7 1347.88 ;
     RECT  1180.7 1325 1180.9 1347.88 ;
     RECT  1179.74 519.86 1181.38 591.88 ;
     RECT  1170.14 1310.72 1181.66 1313.86 ;
     RECT  1180.9 1325 1181.66 1347.46 ;
     RECT  1170.82 610.16 1181.86 610.36 ;
     RECT  1179.94 787.82 1182.82 924.94 ;
     RECT  1178.3 934.4 1183.1 977.86 ;
     RECT  1178.5 1091.06 1183.58 1153.42 ;
     RECT  1173.02 1169.6 1183.58 1210.54 ;
     RECT  1181.66 1308.2 1183.58 1313.86 ;
     RECT  1181.66 1323.32 1183.58 1347.46 ;
     RECT  1181.38 531.2 1183.78 591.88 ;
     RECT  1180.42 1059.98 1183.78 1069.84 ;
     RECT  1159.78 1271.66 1184.06 1276.9 ;
     RECT  1183.78 542.54 1184.74 591.88 ;
     RECT  1184.06 1270.82 1185.22 1276.9 ;
     RECT  1179.94 727.76 1185.5 775 ;
     RECT  1173 -70 1185.98 178 ;
     RECT  1169.18 1219.16 1185.98 1219.78 ;
     RECT  1176.1 1234.28 1185.98 1252.96 ;
     RECT  1185.98 -70 1186.42 179.955 ;
     RECT  1183.1 934.4 1187.42 981.22 ;
     RECT  1183.78 1067.54 1187.42 1069.84 ;
     RECT  1185.98 1219.16 1187.9 1252.96 ;
     RECT  1187.9 1219.16 1188.38 1257.16 ;
     RECT  1188.38 1219.16 1190.78 1262.2 ;
     RECT  1185.22 1270.82 1190.78 1276.48 ;
     RECT  1183.58 1091.06 1191.26 1210.54 ;
     RECT  1190.78 1219.16 1191.26 1276.48 ;
     RECT  1182.62 678.2 1191.74 678.4 ;
     RECT  1180.42 989.84 1191.74 1051.36 ;
     RECT  1175.14 1286.36 1191.74 1299.58 ;
     RECT  1182.82 787.82 1192.22 924.52 ;
     RECT  1160.74 1359.02 1192.22 1359.22 ;
     RECT  1192.22 784.04 1192.7 924.52 ;
     RECT  1187.42 933.14 1192.7 981.22 ;
     RECT  1191.74 989.84 1193.18 1056.82 ;
     RECT  1187.42 1067.54 1193.18 1071.94 ;
     RECT  1183.58 1308.2 1193.18 1347.46 ;
     RECT  1192.22 1359.02 1193.18 1366.78 ;
     RECT  1191.74 677.78 1194.14 678.4 ;
     RECT  1194.14 670.64 1194.62 679.24 ;
     RECT  1191.74 1285.94 1194.62 1299.58 ;
     RECT  1193.18 1308.2 1194.62 1366.78 ;
     RECT  1181.38 519.86 1195.19 520.06 ;
     RECT  1183.78 531.2 1195.19 531.4 ;
     RECT  1184.74 542.54 1195.19 591.46 ;
     RECT  1185.5 647.96 1195.19 648.16 ;
     RECT  1151.14 658.46 1195.19 658.66 ;
     RECT  1194.62 670.64 1195.19 679.66 ;
     RECT  1186.94 696.68 1195.19 696.88 ;
     RECT  1185.5 720.2 1195.19 775 ;
     RECT  1192.7 784.04 1195.19 981.22 ;
     RECT  1193.18 989.84 1195.19 1071.94 ;
     RECT  1159.3 1080.56 1195.19 1080.76 ;
     RECT  1191.26 1091.06 1195.19 1276.48 ;
     RECT  1194.62 1285.94 1195.19 1366.78 ;
     RECT  1195.19 219.14 1200.81 1580.14 ;
     RECT  1200.81 542.54 1201.06 557.86 ;
     RECT  1200.81 709.7 1201.54 774.16 ;
     RECT  1200.81 1170.02 1201.54 1186.18 ;
     RECT  1200.81 1219.16 1201.54 1276.9 ;
     RECT  1200.81 658.46 1202.02 666.22 ;
     RECT  1201.54 717.26 1202.02 774.16 ;
     RECT  1200.81 1308.62 1202.02 1348.3 ;
     RECT  1202.02 1309.46 1202.5 1348.3 ;
     RECT  1200.81 1197.74 1202.98 1208.86 ;
     RECT  1202.5 1337.6 1202.98 1337.8 ;
     RECT  1202.5 1347.26 1202.98 1348.3 ;
     RECT  1201.54 1170.02 1203.46 1176.1 ;
     RECT  1202.98 1197.74 1203.46 1207.6 ;
     RECT  1201.54 1267.88 1203.46 1276.9 ;
     RECT  1202.5 1309.46 1203.46 1321.84 ;
     RECT  1200.81 647.96 1203.94 648.16 ;
     RECT  1201.54 1219.16 1203.94 1256.74 ;
     RECT  1203.46 1312.4 1203.94 1316.38 ;
     RECT  1202.98 1347.26 1203.94 1347.46 ;
     RECT  1200.81 782.78 1204.42 860.68 ;
     RECT  1203.94 1241.42 1204.42 1256.74 ;
     RECT  1200.81 677.78 1204.9 677.98 ;
     RECT  1203.46 1270.82 1204.9 1276.9 ;
     RECT  1204.9 1270.82 1205.38 1276.06 ;
     RECT  1203.94 1313.24 1205.38 1313.44 ;
     RECT  1200.81 1359.02 1205.38 1359.22 ;
     RECT  1202.02 720.2 1205.86 774.16 ;
     RECT  1203.46 1170.86 1205.86 1176.1 ;
     RECT  1201.54 1184.72 1206.34 1186.18 ;
     RECT  1203.46 1207.4 1206.34 1207.6 ;
     RECT  1204.42 835.28 1206.82 860.68 ;
     RECT  1206.34 1185.98 1206.82 1186.18 ;
     RECT  1203.46 1197.74 1206.82 1198.36 ;
     RECT  1200.81 895.34 1207.3 958.96 ;
     RECT  1207.3 909.62 1208.26 958.96 ;
     RECT  1204.42 1241.42 1209.22 1252.96 ;
     RECT  1205.38 1270.82 1209.22 1275.64 ;
     RECT  1200.81 1058.72 1209.5 1082.44 ;
     RECT  1200.81 1091.06 1209.5 1154.26 ;
     RECT  1205.86 722.3 1209.7 774.16 ;
     RECT  1208.26 909.62 1209.7 958.12 ;
     RECT  1209.5 1058.3 1209.7 1154.26 ;
     RECT  1200.81 1286.36 1209.7 1294.96 ;
     RECT  1204.42 783.62 1210.66 822.04 ;
     RECT  1207.3 895.34 1210.66 897.22 ;
     RECT  1209.7 1124.66 1211.62 1154.26 ;
     RECT  1200.81 870.14 1211.9 885.46 ;
     RECT  1211.62 1124.66 1213.06 1128.64 ;
     RECT  1206.82 842 1213.34 860.68 ;
     RECT  1211.9 870.14 1213.34 886.3 ;
     RECT  1200.81 586.64 1214.98 586.84 ;
     RECT  1202.02 658.46 1215.26 658.66 ;
     RECT  1213.34 842 1215.26 886.3 ;
     RECT  1200.81 968.42 1216.7 1048.42 ;
     RECT  1209.7 1058.3 1216.7 1113.94 ;
     RECT  1200.81 568.58 1216.9 568.78 ;
     RECT  1213.06 1124.66 1217.86 1128.22 ;
     RECT  1215.26 652.58 1218.62 658.66 ;
     RECT  1209.7 722.3 1218.62 761.56 ;
     RECT  1218.62 722.3 1220.06 761.98 ;
     RECT  1209.7 773.96 1220.06 774.16 ;
     RECT  1210.66 783.62 1220.54 817.42 ;
     RECT  1215.26 841.16 1220.54 886.3 ;
     RECT  1210.66 897.02 1220.54 897.22 ;
     RECT  1220.06 722.3 1221.22 774.16 ;
     RECT  1205.86 1175.9 1221.22 1176.1 ;
     RECT  1220.54 783.62 1221.7 819.1 ;
     RECT  1209.7 909.62 1221.7 957.7 ;
     RECT  1222.46 632.42 1223.62 632.62 ;
     RECT  1211.62 1137.26 1223.62 1154.26 ;
     RECT  1218.62 652.16 1224.1 658.66 ;
     RECT  1217.86 1128.02 1224.1 1128.22 ;
     RECT  1223.62 1137.26 1224.1 1153.42 ;
     RECT  1216.7 968.42 1225.34 1113.94 ;
     RECT  1224.1 658.46 1226.02 658.66 ;
     RECT  1221.22 755.9 1226.02 774.16 ;
     RECT  1201.06 549.68 1226.5 557.86 ;
     RECT  1223.9 594.2 1226.5 594.4 ;
     RECT  1225.34 968.42 1226.98 1116.88 ;
     RECT  1220.54 833.6 1227.74 897.22 ;
     RECT  1221.7 909.62 1227.74 951.4 ;
     RECT  1226.98 986.48 1228.42 1116.88 ;
     RECT  1227.74 833.6 1228.7 951.4 ;
     RECT  1228.7 831.5 1228.9 951.4 ;
     RECT  1206.82 1198.16 1229.66 1198.36 ;
     RECT  1228.9 831.5 1229.86 950.98 ;
     RECT  1226.98 968.42 1230.14 977.02 ;
     RECT  1230.14 960.44 1230.34 977.02 ;
     RECT  1228.42 986.48 1230.34 1113.94 ;
     RECT  1221.22 722.3 1230.62 747.28 ;
     RECT  1226.5 557.66 1231.3 557.86 ;
     RECT  1230.34 986.48 1232.26 1046.32 ;
     RECT  1229.86 831.5 1232.74 943 ;
     RECT  1230.62 716.84 1233.7 747.28 ;
     RECT  1221.7 783.62 1233.7 818.68 ;
     RECT  1230.14 1332.56 1233.7 1332.76 ;
     RECT  1232.26 986.48 1234.18 1045.9 ;
     RECT  1229.66 1165.82 1234.18 1166.02 ;
     RECT  1233.7 722.3 1234.46 747.28 ;
     RECT  1226.02 756.74 1234.46 774.16 ;
     RECT  1209.22 1241.42 1234.94 1244.98 ;
     RECT  1233.7 783.62 1235.14 797.26 ;
     RECT  1209.5 667.28 1235.42 667.48 ;
     RECT  1234.18 986.48 1235.42 1045.06 ;
     RECT  1209.7 1292.66 1235.42 1294.96 ;
     RECT  1230.34 960.44 1235.62 974.5 ;
     RECT  1235.62 965.06 1236.58 974.5 ;
     RECT  1233.7 806.72 1237.34 818.68 ;
     RECT  1230.34 1056.62 1237.54 1079.08 ;
     RECT  1235.42 659.3 1238.02 667.48 ;
     RECT  1232.74 831.5 1238.3 868.24 ;
     RECT  1230.34 1091.06 1238.3 1113.94 ;
     RECT  1232.74 881.9 1238.78 943 ;
     RECT  1238.3 829.82 1239.74 868.24 ;
     RECT  1235.42 983.96 1239.94 1045.06 ;
     RECT  1238.3 1091.06 1239.94 1121.08 ;
     RECT  1239.94 1091.06 1240.22 1113.94 ;
     RECT  1228.22 1259.48 1240.22 1259.68 ;
     RECT  1209.22 1270.82 1240.22 1271.02 ;
     RECT  1238.02 659.3 1240.42 659.5 ;
     RECT  1240.22 1090.64 1240.42 1113.94 ;
     RECT  1238.78 881.9 1241.66 947.62 ;
     RECT  1235.14 792.02 1241.86 797.26 ;
     RECT  1240.42 1090.64 1242.34 1109.32 ;
     RECT  1224.1 1137.26 1242.34 1143.34 ;
     RECT  1186.42 -70 1243 178 ;
     RECT  1173 1622 1243 1870 ;
     RECT  1237.34 806.72 1243.1 819.1 ;
     RECT  1239.74 829.4 1243.1 868.24 ;
     RECT  1234.46 722.3 1243.3 774.16 ;
     RECT  1239.94 984.38 1243.3 1045.06 ;
     RECT  1242.34 1091.06 1243.3 1109.32 ;
     RECT  1241.66 881.9 1244.06 949.72 ;
     RECT  1243.3 1018.4 1244.26 1038.76 ;
     RECT  1244.26 1018.4 1246.18 1038.34 ;
     RECT  1245.5 1124.24 1246.18 1124.44 ;
     RECT  1243.3 723.98 1246.66 774.16 ;
     RECT  1237.54 1061.66 1246.66 1075.3 ;
     RECT  1243.1 806.72 1246.94 868.24 ;
     RECT  1244.06 881.9 1247.42 950.98 ;
     RECT  1246.18 1018.4 1247.62 1019.02 ;
     RECT  1236.58 965.06 1247.9 973.24 ;
     RECT  1241.86 793.28 1248.1 797.26 ;
     RECT  1246.66 1061.66 1248.1 1071.52 ;
     RECT  1246.94 806.72 1248.58 868.66 ;
     RECT  1246.66 727.76 1249.54 774.16 ;
     RECT  1247.62 1018.4 1249.54 1018.6 ;
     RECT  1241.18 655.52 1249.82 655.72 ;
     RECT  1247.42 881.9 1249.82 952.24 ;
     RECT  1247.9 960.86 1249.82 973.24 ;
     RECT  1249.82 881.9 1250.78 973.24 ;
     RECT  1249.82 655.52 1250.98 656.14 ;
     RECT  1244.54 595.04 1251.46 595.24 ;
     RECT  1248.58 806.72 1251.46 826.66 ;
     RECT  1250.98 655.94 1251.94 656.14 ;
     RECT  1250.78 881.9 1252.22 974.92 ;
     RECT  1243.3 984.38 1252.22 1004.74 ;
     RECT  1239.26 1188.5 1252.7 1188.7 ;
     RECT  1229.66 1198.16 1252.7 1199.2 ;
     RECT  1252.22 881.9 1252.9 1004.74 ;
     RECT  1243.3 1091.06 1253.66 1105.96 ;
     RECT  1233.98 689.54 1253.86 689.74 ;
     RECT  1248.1 795.8 1254.34 797.26 ;
     RECT  1253.66 1090.64 1254.34 1105.96 ;
     RECT  1251.46 806.72 1254.62 819.52 ;
     RECT  1254.34 1091.06 1255.3 1105.96 ;
     RECT  1255.3 1101.14 1256.26 1105.96 ;
     RECT  1252.7 1188.5 1256.74 1199.2 ;
     RECT  1254.62 802.94 1257.22 819.52 ;
     RECT  1256.74 1195.22 1257.22 1199.2 ;
     RECT  1248.58 837.38 1257.7 868.66 ;
     RECT  1249.54 727.76 1257.98 761.56 ;
     RECT  1252.9 881.9 1258.18 950.98 ;
     RECT  1257.7 840.32 1258.46 868.66 ;
     RECT  1257.98 727.34 1259.42 761.56 ;
     RECT  1249.54 770.6 1259.42 774.16 ;
     RECT  1259.42 727.34 1260.1 774.16 ;
     RECT  1248.1 1071.32 1260.1 1071.52 ;
     RECT  1257.22 807.56 1260.38 819.52 ;
     RECT  1243 0 1261 178 ;
     RECT  1243 1622 1261 1800 ;
     RECT  1258.18 927.26 1261.06 950.98 ;
     RECT  1246.18 1030.16 1261.82 1038.34 ;
     RECT  1261.06 928.94 1262.3 950.98 ;
     RECT  1252.9 960.02 1262.3 1004.74 ;
     RECT  1224.1 1153.22 1263.26 1153.42 ;
     RECT  1258.18 881.9 1263.46 918.22 ;
     RECT  1260.38 807.56 1264.7 822.88 ;
     RECT  1260.1 727.76 1265.86 774.16 ;
     RECT  1258.46 840.32 1266.34 871.6 ;
     RECT  1257.22 1196.48 1266.34 1199.2 ;
     RECT  1263.26 1151.12 1267.1 1153.42 ;
     RECT  1267.58 515.24 1268.06 515.44 ;
     RECT  1268.06 515.24 1268.26 516.7 ;
     RECT  1256.26 1105.76 1269.02 1105.96 ;
     RECT  1266.34 847.04 1269.7 871.6 ;
     RECT  1267.1 1151.12 1271.14 1161.82 ;
     RECT  1234.94 1238.48 1271.14 1244.98 ;
     RECT  1259.9 792.44 1271.42 792.64 ;
     RECT  1265.86 773.12 1271.62 774.16 ;
     RECT  1271.42 783.62 1271.9 792.64 ;
     RECT  1264.7 807.56 1271.9 826.66 ;
     RECT  1263.46 882.74 1271.9 918.22 ;
     RECT  1240.22 1259.48 1271.9 1271.02 ;
     RECT  1271.9 882.74 1272.1 919.9 ;
     RECT  1272.1 901.64 1272.86 919.9 ;
     RECT  1262.3 928.94 1272.86 1004.74 ;
     RECT  1235.42 1292.24 1273.82 1294.96 ;
     RECT  1271.9 1259.48 1274.5 1275.22 ;
     RECT  1271.9 783.62 1274.78 826.66 ;
     RECT  1270.94 835.28 1274.78 835.48 ;
     RECT  1255.3 1091.06 1274.98 1091.68 ;
     RECT  1271.14 1153.22 1274.98 1161.82 ;
     RECT  1203.94 1219.16 1275.26 1227.76 ;
     RECT  1274.78 783.62 1276.9 835.48 ;
     RECT  1273.82 1292.24 1277.18 1295.8 ;
     RECT  1275.26 1219.16 1277.38 1229.44 ;
     RECT  1269.7 847.04 1277.86 868.66 ;
     RECT  1277.86 860.48 1278.14 868.66 ;
     RECT  1272.1 882.74 1278.14 890.08 ;
     RECT  1271.14 1241.42 1278.14 1244.98 ;
     RECT  1276.9 783.62 1278.34 826.66 ;
     RECT  1277.38 1219.16 1278.34 1227.76 ;
     RECT  1261.82 1025.96 1280.26 1038.34 ;
     RECT  1272.86 901.64 1280.54 1004.74 ;
     RECT  1269.02 1105.76 1281.22 1113.1 ;
     RECT  1265.86 727.76 1281.7 761.98 ;
     RECT  1262.78 538.76 1282.94 538.96 ;
     RECT  1268.54 548.84 1282.94 549.04 ;
     RECT  1281.7 734.9 1282.94 761.98 ;
     RECT  1271.62 773.96 1282.94 774.16 ;
     RECT  1278.14 860.48 1282.94 890.08 ;
     RECT  1242.34 1137.26 1283.42 1139.98 ;
     RECT  1282.94 860.48 1284.38 893.02 ;
     RECT  1280.54 901.64 1284.38 1010.2 ;
     RECT  1284.38 578.24 1284.86 578.44 ;
     RECT  1278.34 798.74 1285.34 826.66 ;
     RECT  1276.9 835.28 1285.34 835.48 ;
     RECT  1282.94 734.9 1285.54 762.4 ;
     RECT  1285.34 798.74 1286.3 835.48 ;
     RECT  1277.86 847.04 1286.3 848.08 ;
     RECT  1278.34 783.62 1286.78 784.24 ;
     RECT  1283.42 1137.26 1286.98 1143.34 ;
     RECT  1284.38 860.48 1288.7 1010.2 ;
     RECT  1288.7 859.64 1288.9 1010.2 ;
     RECT  1286.78 783.62 1289.18 787.18 ;
     RECT  1271.9 1173.8 1289.66 1174 ;
     RECT  1285.54 736.16 1290.62 762.4 ;
     RECT  1282.94 772.28 1290.62 774.16 ;
     RECT  1281.22 1105.76 1290.82 1109.74 ;
     RECT  1274.98 1153.22 1291.58 1153.42 ;
     RECT  1291.58 1153.22 1291.78 1159.3 ;
     RECT  1260.86 440.48 1292.54 440.68 ;
     RECT  1282.94 538.76 1292.74 549.04 ;
     RECT  1277.18 1286.78 1293.22 1295.8 ;
     RECT  1278.34 1227.56 1293.98 1227.76 ;
     RECT  1278.14 1241.42 1293.98 1248.76 ;
     RECT  1288.9 859.64 1294.18 874.96 ;
     RECT  1289.66 1173.38 1294.66 1174 ;
     RECT  1248.1 1061.66 1294.94 1061.86 ;
     RECT  1286.98 1139.78 1294.94 1143.34 ;
     RECT  1291.78 1153.22 1294.94 1158.88 ;
     RECT  1290.62 736.16 1295.62 774.16 ;
     RECT  1288.9 885.26 1296.1 1010.2 ;
     RECT  1296.1 918.02 1296.58 1010.2 ;
     RECT  1294.18 862.16 1297.82 874.96 ;
     RECT  1292.54 440.48 1298.02 447.82 ;
     RECT  1296.1 885.26 1298.02 909.4 ;
     RECT  1296.58 926.84 1298.02 1010.2 ;
     RECT  1294.94 1139.78 1298.02 1158.88 ;
     RECT  1284.86 578.24 1298.98 580.12 ;
     RECT  1289.18 783.62 1298.98 789.7 ;
     RECT  1293.98 1227.56 1298.98 1248.76 ;
     RECT  1293.5 727.34 1299.26 727.54 ;
     RECT  1295.62 736.16 1299.26 769.12 ;
     RECT  1298.02 447.62 1299.46 447.82 ;
     RECT  1298.02 1139.78 1299.46 1153.42 ;
     RECT  1298.98 783.62 1299.74 787.18 ;
     RECT  1296.38 708.86 1299.94 709.06 ;
     RECT  1299.74 782.78 1300.42 787.18 ;
     RECT  1286.3 798.74 1300.7 849.34 ;
     RECT  1300.22 716 1300.9 716.2 ;
     RECT  1300.7 795.8 1300.9 849.34 ;
     RECT  1298.02 926.84 1301.38 945.1 ;
     RECT  1292.74 538.76 1301.66 538.96 ;
     RECT  1299.74 1123.82 1301.86 1124.02 ;
     RECT  1292.74 548.84 1302.62 549.04 ;
     RECT  1293.22 1286.78 1302.82 1294.96 ;
     RECT  1302.14 639.98 1303.1 640.18 ;
     RECT  1266.34 1199 1303.1 1199.2 ;
     RECT  1298.98 1241.42 1303.58 1248.76 ;
     RECT  1299.46 1151.12 1304.26 1153.42 ;
     RECT  1300.42 782.78 1304.74 784.24 ;
     RECT  1300.9 804.62 1305.22 841.78 ;
     RECT  1300.7 1309.46 1305.22 1309.66 ;
     RECT  1304.74 784.04 1305.7 784.24 ;
     RECT  1300.9 795.8 1306.18 796 ;
     RECT  1274.98 1091.06 1306.66 1091.26 ;
     RECT  1298.02 885.26 1307.42 908.98 ;
     RECT  1296.58 918.02 1307.42 918.22 ;
     RECT  1301.66 538.34 1307.62 538.96 ;
     RECT  1297.82 1211.18 1307.62 1211.38 ;
     RECT  1299.26 727.34 1308.58 769.12 ;
     RECT  1294.66 1173.38 1309.06 1173.58 ;
     RECT  1298.98 1227.56 1309.34 1227.76 ;
     RECT  1303.58 1241.42 1309.34 1249.18 ;
     RECT  1308.58 736.16 1310.02 769.12 ;
     RECT  1302.62 548.84 1310.3 553.24 ;
     RECT  1297.82 862.16 1310.3 876.22 ;
     RECT  1303.1 1195.64 1310.3 1199.2 ;
     RECT  1298.98 578.24 1310.5 578.44 ;
     RECT  1310.02 742.88 1310.5 769.12 ;
     RECT  1305.22 804.62 1310.5 830.44 ;
     RECT  1305.22 841.58 1310.5 841.78 ;
     RECT  1310.3 856.28 1310.5 876.22 ;
     RECT  1298.02 954.56 1310.5 1010.2 ;
     RECT  1309.34 1227.56 1310.5 1249.18 ;
     RECT  1307.42 885.26 1310.78 918.22 ;
     RECT  1301.38 932.72 1310.98 945.1 ;
     RECT  1280.26 1025.96 1311.74 1037.08 ;
     RECT  1310.5 1241.42 1312.22 1249.18 ;
     RECT  1274.5 1259.48 1312.22 1271.02 ;
     RECT  1309.34 519.44 1312.42 519.64 ;
     RECT  1299.46 1139.78 1312.42 1139.98 ;
     RECT  1311.26 655.94 1312.7 656.14 ;
     RECT  1310.5 856.28 1313.66 870.76 ;
     RECT  1310.3 1195.64 1313.86 1205.08 ;
     RECT  1310.98 935.24 1314.14 945.1 ;
     RECT  1310.5 954.56 1314.14 974.08 ;
     RECT  1310.78 882.32 1314.34 918.22 ;
     RECT  1313.66 849.56 1315.3 870.76 ;
     RECT  1261 -70 1315.58 178 ;
     RECT  1314.62 1162.04 1315.58 1162.24 ;
     RECT  1314.34 882.32 1315.78 896.8 ;
     RECT  1310.5 989.84 1315.78 1010.2 ;
     RECT  1315.58 -70 1316.02 179.955 ;
     RECT  1314.14 935.24 1316.26 974.08 ;
     RECT  1311.74 1218.74 1316.26 1218.94 ;
     RECT  1314.62 723.56 1317.22 723.76 ;
     RECT  1314.34 905.42 1317.22 918.22 ;
     RECT  1312.7 655.52 1317.5 656.14 ;
     RECT  1304.26 1153.22 1317.5 1153.42 ;
     RECT  1317.5 1279.64 1318.18 1279.84 ;
     RECT  1315.58 1162.04 1318.46 1166.44 ;
     RECT  1310.3 548.84 1318.94 559.12 ;
     RECT  1310.5 742.88 1318.94 751.06 ;
     RECT  1310.5 761.36 1318.94 769.12 ;
     RECT  1318.94 742.88 1319.14 776.68 ;
     RECT  1316.26 953.72 1319.14 974.08 ;
     RECT  1310.3 592.52 1319.9 592.72 ;
     RECT  1317.5 602.6 1319.9 602.8 ;
     RECT  1319.9 592.52 1320.38 602.8 ;
     RECT  1303.1 639.98 1320.38 640.6 ;
     RECT  1317.5 651.74 1320.38 656.14 ;
     RECT  1316.26 935.24 1321.06 943.42 ;
     RECT  1316.54 704.66 1321.82 704.86 ;
     RECT  1319.14 742.88 1321.82 767.02 ;
     RECT  1310.5 805.88 1321.82 830.44 ;
     RECT  1318.94 548.84 1322.02 566.26 ;
     RECT  1321.82 738.68 1322.3 767.02 ;
     RECT  1315.78 996.98 1322.3 1010.2 ;
     RECT  1321.06 935.24 1322.78 935.44 ;
     RECT  1312.22 1241.42 1322.78 1271.02 ;
     RECT  1256.54 489.2 1323.26 489.4 ;
     RECT  1319.14 776.48 1323.26 776.68 ;
     RECT  1321.82 803.36 1323.26 830.44 ;
     RECT  1322.3 737 1324.22 767.02 ;
     RECT  1315.3 856.28 1324.22 870.76 ;
     RECT  1315.78 884 1324.22 896.8 ;
     RECT  1317.5 1179.68 1324.7 1179.88 ;
     RECT  1322.3 674.84 1325.18 675.04 ;
     RECT  1313.86 1199 1325.18 1205.08 ;
     RECT  1323.74 456.44 1325.66 456.64 ;
     RECT  1321.82 1075.1 1325.66 1075.3 ;
     RECT  1324.22 1086.44 1325.66 1086.64 ;
     RECT  1317.22 908.78 1326.62 918.22 ;
     RECT  1319.14 953.72 1326.62 972.82 ;
     RECT  1311.74 618.14 1327.58 618.34 ;
     RECT  1325.18 674.84 1328.06 676.72 ;
     RECT  1322.3 1124.24 1328.06 1124.44 ;
     RECT  1325.66 455.6 1329.02 456.64 ;
     RECT  1322.3 629.06 1329.5 629.26 ;
     RECT  1320.38 639.98 1329.5 656.14 ;
     RECT  1323.26 799.16 1329.5 830.44 ;
     RECT  1323.26 489.2 1329.98 493.6 ;
     RECT  1322.78 928.52 1329.98 935.44 ;
     RECT  1326.62 946.16 1329.98 972.82 ;
     RECT  1328.06 1121.3 1329.98 1124.44 ;
     RECT  1328.06 569 1330.46 572.98 ;
     RECT  1320.38 591.26 1330.46 602.8 ;
     RECT  1317.5 1151.12 1330.46 1153.42 ;
     RECT  1316.02 -70 1331 178 ;
     RECT  1261 1622 1331 1870 ;
     RECT  1306.46 224.6 1331.19 224.8 ;
     RECT  1329.02 450.56 1331.19 456.64 ;
     RECT  1323.26 474.08 1331.19 474.28 ;
     RECT  1329.98 489.2 1331.19 497.38 ;
     RECT  1326.62 506 1331.19 506.2 ;
     RECT  1322.3 526.58 1331.19 526.78 ;
     RECT  1307.62 538.34 1331.19 538.54 ;
     RECT  1322.02 548.84 1331.19 559.12 ;
     RECT  1330.46 569 1331.19 580.96 ;
     RECT  1330.46 591.26 1331.19 606.58 ;
     RECT  1327.58 617.72 1331.19 618.34 ;
     RECT  1329.5 629.06 1331.19 656.14 ;
     RECT  1330.94 664.76 1331.19 664.96 ;
     RECT  1328.06 674.84 1331.19 683.44 ;
     RECT  1321.82 697.1 1331.19 704.86 ;
     RECT  1324.22 735.32 1331.19 767.02 ;
     RECT  1323.26 776.48 1331.19 777.1 ;
     RECT  1329.5 795.8 1331.19 833.8 ;
     RECT  1324.22 856.28 1331.19 896.8 ;
     RECT  1326.62 905.42 1331.19 918.22 ;
     RECT  1329.98 928.52 1331.19 972.82 ;
     RECT  1322.3 996.98 1331.19 1010.62 ;
     RECT  1311.74 1025.96 1331.19 1045.48 ;
     RECT  1294.94 1054.94 1331.19 1061.86 ;
     RECT  1325.66 1075.1 1331.19 1086.64 ;
     RECT  1290.82 1105.76 1331.19 1105.96 ;
     RECT  1329.98 1121.3 1331.19 1128.22 ;
     RECT  1330.46 1150.7 1331.19 1153.42 ;
     RECT  1318.46 1162.04 1331.19 1166.86 ;
     RECT  1324.7 1179.68 1331.19 1182.82 ;
     RECT  1325.18 1199 1331.19 1206.76 ;
     RECT  1310.5 1227.56 1331.19 1228.18 ;
     RECT  1322.78 1241.42 1331.19 1271.44 ;
     RECT  1302.82 1292.24 1331.19 1294.96 ;
     RECT  1326.14 1317.44 1331.19 1317.64 ;
     RECT  1331.19 215.36 1336.81 1583.92 ;
     RECT  1336.81 1124.24 1336.9 1128.64 ;
     RECT  1336.81 489.2 1337.38 559.12 ;
     RECT  1336.81 664.76 1337.38 683.44 ;
     RECT  1336.81 1199 1337.38 1227.76 ;
     RECT  1336.81 1236.8 1337.38 1275.64 ;
     RECT  1336.81 605.96 1337.86 620.02 ;
     RECT  1336.81 1086.44 1337.86 1113.1 ;
     RECT  1336.81 1288.04 1337.86 1295.38 ;
     RECT  1336.81 742.88 1338.34 781.72 ;
     RECT  1336.81 885.26 1338.34 972.82 ;
     RECT  1337.86 1091.48 1338.34 1113.1 ;
     RECT  1337.38 1236.8 1338.34 1271.44 ;
     RECT  1336.81 568.16 1338.82 591.46 ;
     RECT  1336.81 856.28 1338.82 874.96 ;
     RECT  1338.34 905.84 1338.82 972.82 ;
     RECT  1336.9 1128.44 1338.82 1128.64 ;
     RECT  1338.34 1241 1338.82 1271.44 ;
     RECT  1337.86 1290.14 1338.82 1295.38 ;
     RECT  1337.38 500.96 1339.3 511.66 ;
     RECT  1337.38 527 1339.3 559.12 ;
     RECT  1338.82 568.58 1339.3 591.46 ;
     RECT  1337.86 606.38 1339.3 620.02 ;
     RECT  1336.81 790.76 1339.3 822.04 ;
     RECT  1336.81 832.34 1339.3 836.32 ;
     RECT  1336.81 1073 1339.3 1075.3 ;
     RECT  1338.34 1101.56 1339.3 1113.1 ;
     RECT  1337.38 1215.8 1339.3 1227.76 ;
     RECT  1338.82 1241 1339.3 1245.4 ;
     RECT  1338.82 1254.44 1339.3 1271.44 ;
     RECT  1339.3 527 1339.78 534.76 ;
     RECT  1338.34 742.88 1339.78 751.48 ;
     RECT  1338.82 905.84 1339.78 912.76 ;
     RECT  1339.3 1222.52 1339.78 1227.76 ;
     RECT  1339.3 568.58 1340.26 572.98 ;
     RECT  1339.3 791.6 1340.26 822.04 ;
     RECT  1338.82 856.28 1340.26 864.88 ;
     RECT  1336.81 474.08 1340.74 478.48 ;
     RECT  1336.81 629.06 1340.74 656.14 ;
     RECT  1336.81 697.1 1340.74 705.28 ;
     RECT  1340.26 799.16 1340.74 799.36 ;
     RECT  1338.82 923.9 1340.74 972.82 ;
     RECT  1340.74 629.06 1341.22 633.46 ;
     RECT  1339.3 606.38 1341.7 617.92 ;
     RECT  1340.26 856.28 1341.7 864.04 ;
     RECT  1340.74 928.52 1341.7 972.82 ;
     RECT  1337.38 1199 1341.7 1205.08 ;
     RECT  1336.81 450.56 1342.18 464.2 ;
     RECT  1341.7 928.52 1342.18 964.42 ;
     RECT  1339.78 1224.62 1342.18 1227.76 ;
     RECT  1342.18 450.56 1342.66 457.9 ;
     RECT  1339.78 746.24 1344.1 751.48 ;
     RECT  1339.3 1075.1 1344.1 1075.3 ;
     RECT  1339.3 548.84 1344.58 559.12 ;
     RECT  1340.26 807.98 1344.58 822.04 ;
     RECT  1341.7 863.42 1345.54 864.04 ;
     RECT  1342.18 964.22 1345.54 964.42 ;
     RECT  1338.34 766.82 1346.02 777.1 ;
     RECT  1338.82 873.92 1346.02 874.96 ;
     RECT  1336.81 1025.96 1346.02 1037.08 ;
     RECT  1344.58 818.9 1346.5 822.04 ;
     RECT  1338.34 885.26 1346.78 890.5 ;
     RECT  1336.81 1309.88 1346.78 1321 ;
     RECT  1342.18 928.52 1346.98 953.5 ;
     RECT  1346.78 885.26 1347.46 897.64 ;
     RECT  1346.98 928.52 1347.94 942.16 ;
     RECT  1346.78 1306.52 1347.94 1321 ;
     RECT  1340.74 644.18 1348.42 656.14 ;
     RECT  1339.3 1241.42 1348.7 1245.4 ;
     RECT  1339.3 1256.96 1348.9 1271.44 ;
     RECT  1331 0 1349 178 ;
     RECT  1331 1622 1349 1800 ;
     RECT  1339.3 584.96 1349.18 591.46 ;
     RECT  1337.38 664.76 1349.18 664.96 ;
     RECT  1337.38 675.26 1349.18 683.44 ;
     RECT  1339.78 531.62 1349.38 534.76 ;
     RECT  1340.74 697.1 1349.66 704.86 ;
     RECT  1347.46 885.26 1350.14 890.5 ;
     RECT  1345.54 863.42 1350.34 863.62 ;
     RECT  1349.66 697.1 1350.82 705.28 ;
     RECT  1346.02 874.76 1351.1 874.96 ;
     RECT  1350.14 883.58 1351.1 890.5 ;
     RECT  1351.1 874.76 1351.3 890.5 ;
     RECT  1339.78 912.56 1351.3 912.76 ;
     RECT  1336.81 988.58 1351.3 1010.2 ;
     RECT  1339.3 1105.76 1351.3 1113.1 ;
     RECT  1350.82 700.04 1352.26 705.28 ;
     RECT  1340.74 474.08 1352.74 474.28 ;
     RECT  1342.66 450.56 1353.7 456.64 ;
     RECT  1341.22 633.26 1353.7 633.46 ;
     RECT  1350.14 849.14 1353.7 849.34 ;
     RECT  1351.3 881.06 1353.7 890.5 ;
     RECT  1340.26 572.78 1353.98 572.98 ;
     RECT  1353.98 572.78 1354.18 574.66 ;
     RECT  1339.3 832.34 1354.18 833.8 ;
     RECT  1353.7 881.06 1354.66 886.3 ;
     RECT  1353.7 450.56 1354.94 453.28 ;
     RECT  1354.18 574.46 1355.14 574.66 ;
     RECT  1346.98 953.3 1355.14 953.5 ;
     RECT  1347.94 1317.44 1355.14 1321 ;
     RECT  1353.02 783.62 1355.42 783.82 ;
     RECT  1346.5 821.84 1355.62 822.04 ;
     RECT  1354.66 883.16 1355.62 886.3 ;
     RECT  1349.18 583.28 1355.9 591.46 ;
     RECT  1344.58 807.98 1355.9 808.18 ;
     RECT  1349.18 664.76 1356.1 683.44 ;
     RECT  1346.02 766.82 1356.1 773.74 ;
     RECT  1341.7 606.38 1356.58 610.78 ;
     RECT  1355.9 806.72 1356.58 808.18 ;
     RECT  1348.42 644.18 1357.06 651.94 ;
     RECT  1344.1 746.66 1357.06 751.48 ;
     RECT  1347.94 941.96 1357.06 942.16 ;
     RECT  1336.81 1162.04 1357.06 1182.82 ;
     RECT  1355.9 583.28 1357.34 593.98 ;
     RECT  1342.18 1227.56 1357.34 1227.76 ;
     RECT  1357.34 581.18 1357.54 593.98 ;
     RECT  1356.58 606.38 1357.54 606.58 ;
     RECT  1355.42 783.62 1357.54 784.24 ;
     RECT  1355.62 883.16 1357.54 885.46 ;
     RECT  1357.06 1173.38 1357.54 1182.82 ;
     RECT  1356.1 664.76 1357.82 683.02 ;
     RECT  1357.54 593.78 1358.02 593.98 ;
     RECT  1356.1 766.82 1358.02 768.7 ;
     RECT  1354.18 833.6 1358.02 833.8 ;
     RECT  1357.54 883.58 1358.02 885.46 ;
     RECT  1357.06 747.92 1358.3 751.48 ;
     RECT  1356.38 977.24 1358.3 977.44 ;
     RECT  1348.7 1241.42 1358.3 1245.82 ;
     RECT  1348.9 1256.96 1358.3 1271.02 ;
     RECT  1336.81 224.6 1358.5 224.8 ;
     RECT  1357.54 581.18 1358.5 585.16 ;
     RECT  1358.3 747.92 1358.5 758.2 ;
     RECT  1357.54 783.62 1358.5 783.82 ;
     RECT  1357.34 1227.56 1358.5 1228.6 ;
     RECT  1338.82 1292.24 1358.5 1295.38 ;
     RECT  1352.26 704.24 1358.78 705.28 ;
     RECT  1356.58 806.72 1358.98 806.92 ;
     RECT  1357.54 1173.38 1359.46 1179.88 ;
     RECT  1357.06 1162.04 1359.94 1163.92 ;
     RECT  1344.58 550.1 1360.42 559.12 ;
     RECT  1355.42 440.06 1360.7 440.26 ;
     RECT  1357.82 663.5 1360.7 683.02 ;
     RECT  1339.3 506 1360.9 511.66 ;
     RECT  1360.7 662.24 1360.9 683.02 ;
     RECT  1358.5 758 1360.9 758.2 ;
     RECT  1358.02 768.5 1360.9 768.7 ;
     RECT  1359.46 1178 1360.9 1179.88 ;
     RECT  1358.3 977.24 1361.18 979.54 ;
     RECT  1358.78 704.24 1361.38 708.64 ;
     RECT  1341.7 1199 1362.14 1199.2 ;
     RECT  1362.14 855.44 1362.62 855.64 ;
     RECT  1346.02 1025.96 1362.62 1030.36 ;
     RECT  1336.81 1054.94 1362.62 1061.86 ;
     RECT  1362.14 1199 1362.82 1205.5 ;
     RECT  1360.9 662.24 1363.1 662.44 ;
     RECT  1358.3 1241.42 1363.1 1271.02 ;
     RECT  1361.18 977.24 1363.58 982.48 ;
     RECT  1362.62 855.44 1363.78 863.62 ;
     RECT  1358.3 1324.58 1363.78 1324.78 ;
     RECT  1360.7 842 1364.26 842.2 ;
     RECT  1363.78 855.44 1364.26 855.64 ;
     RECT  1351.3 996.98 1364.54 1010.2 ;
     RECT  1358.5 1227.56 1364.54 1227.76 ;
     RECT  1360.7 439.22 1364.74 440.26 ;
     RECT  1363.1 1236.8 1364.74 1271.02 ;
     RECT  1360.7 1282.16 1365.5 1282.36 ;
     RECT  1358.5 1292.24 1365.5 1294.96 ;
     RECT  1347.94 1306.52 1365.7 1306.72 ;
     RECT  1362.62 1025.96 1365.98 1037.92 ;
     RECT  1365.5 1093.16 1366.18 1093.36 ;
     RECT  1365.98 1025.96 1366.46 1041.28 ;
     RECT  1336.81 1151.12 1366.46 1153.42 ;
     RECT  1359.94 1162.04 1366.46 1162.24 ;
     RECT  1351.3 1105.76 1366.94 1105.96 ;
     RECT  1366.46 1025.96 1367.42 1041.7 ;
     RECT  1365.98 562.28 1367.62 562.48 ;
     RECT  1363.1 654.26 1367.62 662.44 ;
     RECT  1367.62 659.72 1368.1 662.44 ;
     RECT  1360.7 620.66 1368.38 627.16 ;
     RECT  1366.94 1105.76 1368.38 1109.74 ;
     RECT  1364.54 992.78 1368.58 1010.2 ;
     RECT  1363.58 977.24 1368.86 984.16 ;
     RECT  1368.58 992.78 1368.86 1002.22 ;
     RECT  1366.46 1151.12 1368.86 1162.24 ;
     RECT  1368.38 617.3 1369.34 627.16 ;
     RECT  1364.74 440.06 1369.54 440.26 ;
     RECT  1368.86 1151.12 1369.82 1169.8 ;
     RECT  1368.1 659.72 1370.5 659.92 ;
     RECT  1367.42 1018.82 1370.5 1041.7 ;
     RECT  1368.38 1105.76 1370.5 1117.72 ;
     RECT  1357.06 644.18 1370.78 644.38 ;
     RECT  1362.62 1054.94 1370.78 1067.74 ;
     RECT  1367.9 1128.44 1370.78 1128.64 ;
     RECT  1369.82 1151.12 1370.78 1173.58 ;
     RECT  1349.38 531.62 1371.26 531.82 ;
     RECT  1370.78 640.4 1371.26 644.38 ;
     RECT  1360.9 511.46 1371.46 511.66 ;
     RECT  1370.5 1038.56 1371.74 1041.7 ;
     RECT  1365.5 1282.16 1371.74 1294.96 ;
     RECT  1362.14 1083.08 1371.94 1083.28 ;
     RECT  1370.78 1149.44 1371.94 1173.58 ;
     RECT  1364.54 1219.16 1372.22 1227.76 ;
     RECT  1364.74 1241.42 1372.22 1271.02 ;
     RECT  1371.74 1280.06 1372.22 1294.96 ;
     RECT  1369.34 613.94 1372.9 627.16 ;
     RECT  1370.5 1105.76 1373.86 1109.74 ;
     RECT  1358.5 747.92 1374.62 748.12 ;
     RECT  1354.94 448.88 1375.1 453.28 ;
     RECT  1358.5 584.96 1375.1 585.16 ;
     RECT  1361.38 704.24 1375.1 704.44 ;
     RECT  1375.1 584.12 1375.3 585.16 ;
     RECT  1370.78 1052.84 1375.58 1067.74 ;
     RECT  1373.86 1105.76 1375.58 1105.96 ;
     RECT  1362.82 1199 1375.58 1199.2 ;
     RECT  1372.22 1215.38 1375.58 1227.76 ;
     RECT  1372.22 1241.42 1375.58 1294.96 ;
     RECT  1360.42 550.1 1376.06 550.3 ;
     RECT  1375.1 704.24 1376.06 711.58 ;
     RECT  1375.58 1052.84 1376.06 1068.16 ;
     RECT  1371.74 1038.56 1376.26 1042.54 ;
     RECT  1371.26 530.78 1376.54 531.82 ;
     RECT  1371.26 636.62 1376.54 644.38 ;
     RECT  1376.06 704.24 1376.54 715.78 ;
     RECT  1347.94 928.52 1376.54 928.72 ;
     RECT  1371.94 1153.22 1376.54 1173.58 ;
     RECT  1375.58 1215.38 1377.02 1294.96 ;
     RECT  1375.3 584.12 1377.22 584.32 ;
     RECT  1373.66 894.08 1377.22 902.26 ;
     RECT  1376.54 530.78 1377.5 535.18 ;
     RECT  1376.06 1052.84 1377.5 1075.72 ;
     RECT  1376.54 702.56 1377.7 715.78 ;
     RECT  1376.26 1038.56 1377.7 1038.76 ;
     RECT  1377.5 1051.58 1377.98 1075.72 ;
     RECT  1377.02 1211.18 1377.98 1294.96 ;
     RECT  1377.98 1210.76 1378.18 1294.96 ;
     RECT  1368.86 977.24 1378.46 1002.22 ;
     RECT  1377.5 525.32 1378.66 535.18 ;
     RECT  1377.5 874.76 1378.94 874.96 ;
     RECT  1358.02 885.26 1378.94 885.46 ;
     RECT  1375.58 1100.3 1378.94 1105.96 ;
     RECT  1378.18 1290.98 1379.14 1294.96 ;
     RECT  1376.54 1153.22 1379.62 1174 ;
     RECT  1376.54 927.26 1379.9 928.72 ;
     RECT  1375.1 758 1380.38 758.2 ;
     RECT  1378.94 874.76 1380.38 885.46 ;
     RECT  1378.46 977.24 1380.38 1003.06 ;
     RECT  1375.58 1193.54 1380.38 1199.2 ;
     RECT  1380.38 758 1380.58 763.24 ;
     RECT  1379.9 924.74 1380.58 928.72 ;
     RECT  1380.38 977.24 1380.58 1007.68 ;
     RECT  1369.34 1313.24 1380.58 1313.44 ;
     RECT  1374.62 863.84 1380.86 864.04 ;
     RECT  1380.38 874.34 1380.86 885.46 ;
     RECT  1377.98 1048.64 1381.54 1075.72 ;
     RECT  1379.14 1292.24 1381.82 1294.96 ;
     RECT  1380.58 977.24 1382.02 982.48 ;
     RECT  1380.58 927.26 1382.5 928.72 ;
     RECT  1378.18 1210.76 1382.5 1277.32 ;
     RECT  1376.54 632.42 1382.98 644.38 ;
     RECT  1378.94 1094 1382.98 1105.96 ;
     RECT  1377.22 897.44 1383.26 902.26 ;
     RECT  1382.98 632.84 1383.74 644.38 ;
     RECT  1383.74 632.84 1384.22 648.58 ;
     RECT  1381.54 1048.64 1384.42 1051.78 ;
     RECT  1380.86 860.06 1384.9 885.46 ;
     RECT  1370.5 1018.82 1385.18 1026.58 ;
     RECT  1375.1 965.06 1386.14 965.26 ;
     RECT  1383.26 897.44 1387.3 909.4 ;
     RECT  1384.9 867.2 1387.78 885.46 ;
     RECT  1386.62 802.94 1388.54 803.14 ;
     RECT  1381.54 1061.66 1389.22 1075.72 ;
     RECT  1379.62 1158.68 1389.22 1174 ;
     RECT  1374.62 741.2 1389.7 748.12 ;
     RECT  1382.98 1097.78 1389.7 1105.96 ;
     RECT  1377.7 702.56 1389.98 704.44 ;
     RECT  1377.7 715.58 1389.98 715.78 ;
     RECT  1380.58 992.78 1389.98 1007.68 ;
     RECT  1360.9 672.32 1390.46 683.02 ;
     RECT  1381.82 1292.24 1390.46 1302.52 ;
     RECT  1387.58 788.24 1390.94 788.44 ;
     RECT  1389.98 992.36 1390.94 1007.68 ;
     RECT  1382.02 977.24 1391.42 979.54 ;
     RECT  1390.94 988.58 1391.42 1007.68 ;
     RECT  1389.7 746.24 1391.9 748.12 ;
     RECT  1382.5 928.52 1391.9 928.72 ;
     RECT  1391.42 436.7 1392.38 436.9 ;
     RECT  1375.1 448.04 1392.38 453.28 ;
     RECT  1389.98 702.56 1392.86 715.78 ;
     RECT  1386.62 954.14 1392.86 954.34 ;
     RECT  1386.14 965.06 1392.86 965.68 ;
     RECT  1385.18 1017.98 1392.86 1026.58 ;
     RECT  1370.78 1122.98 1392.86 1128.64 ;
     RECT  1387.78 874.34 1393.82 885.46 ;
     RECT  1385.66 602.6 1394.3 602.8 ;
     RECT  1391.9 920.12 1394.3 928.72 ;
     RECT  1389.22 1172.96 1394.78 1174 ;
     RECT  1378.66 530.78 1395.26 535.18 ;
     RECT  1390.94 784.04 1395.26 788.44 ;
     RECT  1386.62 512.3 1395.74 512.5 ;
     RECT  1395.26 526.16 1395.74 535.18 ;
     RECT  1391.42 977.24 1395.74 1007.68 ;
     RECT  1389.22 1158.68 1395.74 1162.24 ;
     RECT  1395.74 976.82 1396.22 1007.68 ;
     RECT  1380.38 1193.54 1396.22 1200.46 ;
     RECT  1392.86 1119.62 1396.7 1128.64 ;
     RECT  1386.62 1143.56 1396.7 1143.76 ;
     RECT  1390.46 1290.56 1396.7 1302.52 ;
     RECT  1394.78 586.22 1397.18 586.42 ;
     RECT  1372.9 613.94 1397.18 620.86 ;
     RECT  1384.22 632.84 1397.18 656.98 ;
     RECT  1395.74 1157.42 1397.18 1162.24 ;
     RECT  1396.22 1193.54 1397.18 1201.3 ;
     RECT  1396.7 1290.56 1397.18 1306.72 ;
     RECT  1395.74 512.3 1397.66 535.18 ;
     RECT  1397.18 572.78 1397.66 572.98 ;
     RECT  1392.86 953.72 1397.66 965.68 ;
     RECT  1396.22 976.4 1397.66 1007.68 ;
     RECT  1389.7 1098.2 1397.66 1105.96 ;
     RECT  1396.7 1119.62 1397.66 1143.76 ;
     RECT  1397.18 1290.56 1397.66 1309.66 ;
     RECT  1393.34 941.96 1398.14 942.16 ;
     RECT  1397.66 953.72 1398.14 1007.68 ;
     RECT  1392.86 1017.98 1398.14 1029.94 ;
     RECT  1337.38 489.2 1398.62 489.4 ;
     RECT  1392.86 702.56 1398.62 723.76 ;
     RECT  1398.14 953.72 1398.62 1029.94 ;
     RECT  1394.78 1172.96 1398.62 1177.36 ;
     RECT  1382.5 1211.18 1398.62 1277.32 ;
     RECT  1397.66 1290.56 1398.62 1312.18 ;
     RECT  1376.06 550.1 1399.1 553.24 ;
     RECT  1392.38 436.7 1399.19 453.28 ;
     RECT  1381.34 462.74 1399.19 462.94 ;
     RECT  1398.62 482.9 1399.19 489.4 ;
     RECT  1397.66 512.3 1399.19 536.02 ;
     RECT  1399.1 550.1 1399.19 558.7 ;
     RECT  1397.66 572.78 1399.19 576.34 ;
     RECT  1397.18 586.22 1399.19 590.2 ;
     RECT  1394.3 602.6 1399.19 603.22 ;
     RECT  1397.18 613.94 1399.19 656.98 ;
     RECT  1390.46 666.86 1399.19 683.02 ;
     RECT  1398.62 696.68 1399.19 723.76 ;
     RECT  1391.9 746.24 1399.19 754 ;
     RECT  1380.58 763.04 1399.19 763.24 ;
     RECT  1395.26 780.68 1399.19 788.86 ;
     RECT  1388.54 800 1399.19 803.14 ;
     RECT  1398.62 858.8 1399.19 859 ;
     RECT  1393.82 874.34 1399.19 887.14 ;
     RECT  1387.3 897.44 1399.19 902.26 ;
     RECT  1394.3 916.34 1399.19 928.72 ;
     RECT  1398.14 940.28 1399.19 942.16 ;
     RECT  1398.62 951.62 1399.19 1029.94 ;
     RECT  1384.42 1051.58 1399.19 1051.78 ;
     RECT  1389.22 1061.66 1399.19 1061.86 ;
     RECT  1389.22 1075.52 1399.19 1075.72 ;
     RECT  1397.66 1098.2 1399.19 1143.76 ;
     RECT  1397.18 1154.48 1399.19 1162.24 ;
     RECT  1398.62 1170.86 1399.19 1177.36 ;
     RECT  1397.18 1189.34 1399.19 1201.3 ;
     RECT  1398.62 1211.18 1399.19 1312.18 ;
     RECT  1394.78 1328.36 1399.19 1328.56 ;
     RECT  1349 -70 1403.9 178 ;
     RECT  1399.19 219.14 1404.81 1580.14 ;
     RECT  1404.81 432.92 1405.06 453.7 ;
     RECT  1404.81 780.68 1405.54 803.14 ;
     RECT  1404.81 858.8 1405.54 859 ;
     RECT  1404.81 1120.88 1405.54 1121.08 ;
     RECT  1404.81 1292.24 1405.54 1302.52 ;
     RECT  1404.81 545.06 1406.02 558.7 ;
     RECT  1404.81 590 1406.02 602.8 ;
     RECT  1405.54 784.04 1406.02 803.14 ;
     RECT  1405.06 432.92 1406.5 436.9 ;
     RECT  1404.81 667.7 1406.5 683.02 ;
     RECT  1404.81 696.68 1406.5 719.14 ;
     RECT  1406.02 784.04 1406.5 796.84 ;
     RECT  1404.81 909.2 1406.5 910.24 ;
     RECT  1404.81 953.72 1406.5 1008.94 ;
     RECT  1404.81 1211.18 1406.5 1227.76 ;
     RECT  1403.9 -70 1406.98 179.44 ;
     RECT  1406.5 788.24 1406.98 796.84 ;
     RECT  1404.81 1311.98 1406.98 1312.18 ;
     RECT  1404.81 615.62 1407.46 658.66 ;
     RECT  1406.98 788.24 1407.46 788.86 ;
     RECT  1404.81 1143.56 1407.46 1154.68 ;
     RECT  1406.02 546.32 1407.94 558.7 ;
     RECT  1404.81 577.4 1407.94 577.6 ;
     RECT  1406.5 718.1 1408.42 719.14 ;
     RECT  1404.81 1168.76 1408.42 1199.2 ;
     RECT  1404.81 462.74 1408.9 465.88 ;
     RECT  1404.81 512.3 1408.9 512.5 ;
     RECT  1404.81 1075.52 1408.9 1078.66 ;
     RECT  1407.46 1143.56 1408.9 1151.32 ;
     RECT  1407.46 615.62 1409.38 656.98 ;
     RECT  1408.9 1078.46 1409.38 1078.66 ;
     RECT  1404.81 1098.2 1409.38 1110.16 ;
     RECT  1404.81 737.84 1409.86 738.04 ;
     RECT  1404.81 1018.4 1409.86 1026.58 ;
     RECT  1406.5 696.68 1410.34 704.44 ;
     RECT  1406.5 962.12 1410.34 1008.94 ;
     RECT  1409.38 1099.46 1410.34 1110.16 ;
     RECT  1404.81 746.66 1410.82 748.12 ;
     RECT  1408.42 1168.76 1410.82 1184.08 ;
     RECT  1405.06 448.04 1411.3 453.7 ;
     RECT  1407.94 546.32 1411.3 554.5 ;
     RECT  1406.5 672.32 1411.3 683.02 ;
     RECT  1407.46 788.66 1411.3 788.86 ;
     RECT  1410.34 1008.74 1411.3 1008.94 ;
     RECT  1410.34 1105.76 1411.3 1110.16 ;
     RECT  1410.34 962.12 1411.78 969.46 ;
     RECT  1411.3 546.32 1412.26 546.52 ;
     RECT  1404.81 885.26 1412.74 897.64 ;
     RECT  1408.9 1150.7 1412.74 1151.32 ;
     RECT  1412.74 1151.12 1413.7 1151.32 ;
     RECT  1404.81 489.2 1414.46 489.4 ;
     RECT  1409.38 615.62 1414.66 640.18 ;
     RECT  1408.42 718.1 1414.94 718.3 ;
     RECT  1405.54 1292.24 1415.14 1302.1 ;
     RECT  1406.02 592.1 1415.9 601.12 ;
     RECT  1412.74 885.26 1415.9 887.56 ;
     RECT  1404.81 923.48 1415.9 928.72 ;
     RECT  1409.86 1026.38 1415.9 1026.58 ;
     RECT  1414.66 617.72 1416.1 640.18 ;
     RECT  1416.1 618.14 1417.54 640.18 ;
     RECT  1404.81 1241.42 1417.54 1279.84 ;
     RECT  1412.74 897.44 1418.02 897.64 ;
     RECT  1417.54 1241.42 1418.5 1272.28 ;
     RECT  1415.9 882.74 1418.78 887.56 ;
     RECT  1406.98 -70 1419 178 ;
     RECT  1349 1622 1419 1870 ;
     RECT  1415.9 920.54 1419.74 928.72 ;
     RECT  1410.34 704.24 1420.22 704.44 ;
     RECT  1418.78 874.76 1420.22 887.56 ;
     RECT  1406.5 432.92 1420.42 433.12 ;
     RECT  1418.5 1241.42 1420.7 1271.02 ;
     RECT  1410.34 980.18 1421.18 999.7 ;
     RECT  1418.78 1010.84 1421.18 1011.04 ;
     RECT  1406.5 1211.18 1422.14 1213.06 ;
     RECT  1406.5 1225.46 1422.14 1227.76 ;
     RECT  1420.22 697.52 1422.62 704.44 ;
     RECT  1411.3 1105.76 1423.1 1105.96 ;
     RECT  1418.78 1115.84 1423.1 1116.04 ;
     RECT  1422.14 1211.18 1423.3 1227.76 ;
     RECT  1411.3 675.26 1423.58 683.02 ;
     RECT  1422.62 692.48 1423.58 704.44 ;
     RECT  1420.22 870.98 1423.58 887.56 ;
     RECT  1418.78 783.2 1423.78 783.4 ;
     RECT  1411.78 969.26 1423.78 969.46 ;
     RECT  1414.94 715.58 1424.54 718.3 ;
     RECT  1417.34 957.92 1424.74 958.12 ;
     RECT  1419.74 919.28 1425.5 928.72 ;
     RECT  1417.54 618.14 1425.7 625.48 ;
     RECT  1423.58 675.26 1425.7 704.44 ;
     RECT  1415.9 592.1 1425.98 605.74 ;
     RECT  1415.14 1292.24 1426.46 1300.42 ;
     RECT  1425.5 563.96 1426.66 565 ;
     RECT  1426.46 1136.42 1427.42 1136.62 ;
     RECT  1410.82 1173.8 1427.42 1184.08 ;
     RECT  1423.1 1105.76 1427.9 1116.04 ;
     RECT  1425.7 618.14 1428.1 618.34 ;
     RECT  1423.58 870.98 1428.38 888.4 ;
     RECT  1427.42 1131.38 1428.38 1136.62 ;
     RECT  1409.38 648.8 1428.58 649 ;
     RECT  1428.38 1131.38 1428.58 1137.04 ;
     RECT  1415.9 1026.38 1429.54 1031.62 ;
     RECT  1427.42 1171.28 1429.54 1184.08 ;
     RECT  1423.58 765.56 1429.82 765.76 ;
     RECT  1408.9 465.68 1430.3 465.88 ;
     RECT  1423.3 1211.18 1430.98 1213.06 ;
     RECT  1430.3 822.26 1431.74 822.46 ;
     RECT  1428.86 834.44 1431.74 834.64 ;
     RECT  1424.06 905.42 1431.74 905.62 ;
     RECT  1425.5 915.92 1431.74 928.72 ;
     RECT  1421.18 980.18 1431.94 1011.04 ;
     RECT  1424.54 715.58 1432.22 720.4 ;
     RECT  1429.54 1026.38 1432.22 1026.58 ;
     RECT  1431.94 1002.86 1432.42 1011.04 ;
     RECT  1431.74 905.42 1432.9 928.72 ;
     RECT  1428.38 867.62 1433.38 888.4 ;
     RECT  1426.94 780.26 1433.66 781.3 ;
     RECT  1426.46 799.58 1433.66 799.78 ;
     RECT  1426.46 1292.24 1433.86 1305.88 ;
     RECT  1432.7 849.14 1434.14 849.34 ;
     RECT  1421.18 664.34 1434.34 664.54 ;
     RECT  1432.42 1010.84 1434.34 1011.04 ;
     RECT  1433.38 867.62 1434.82 882.52 ;
     RECT  1431.94 980.18 1435.78 992.56 ;
     RECT  1404.81 526.16 1436.06 531.82 ;
     RECT  1434.82 876.86 1436.26 882.52 ;
     RECT  1423.3 1225.46 1436.54 1227.76 ;
     RECT  1420.7 1240.58 1436.54 1271.02 ;
     RECT  1436.26 876.86 1436.74 877.9 ;
     RECT  1419 0 1437 178 ;
     RECT  1419 1622 1437 1800 ;
     RECT  1431.74 822.26 1437.02 834.64 ;
     RECT  1425.98 584.12 1437.7 607.42 ;
     RECT  1432.9 909.2 1438.66 928.72 ;
     RECT  1432.7 947 1438.66 947.2 ;
     RECT  1433.66 798.32 1438.94 799.78 ;
     RECT  1429.54 1173.8 1438.94 1184.08 ;
     RECT  1408.42 1196.06 1438.94 1199.2 ;
     RECT  1417.54 636.62 1439.42 640.18 ;
     RECT  1438.94 1173.8 1439.42 1199.2 ;
     RECT  1430.98 1211.18 1439.42 1211.8 ;
     RECT  1436.06 519.86 1439.62 531.82 ;
     RECT  1439.42 1173.8 1440.1 1216 ;
     RECT  1436.54 1225.46 1440.1 1271.02 ;
     RECT  1429.82 765.14 1440.38 765.76 ;
     RECT  1433.66 780.26 1440.38 785.08 ;
     RECT  1425.98 739.1 1440.58 739.3 ;
     RECT  1438.94 795.38 1440.58 799.78 ;
     RECT  1436.74 877.7 1440.58 877.9 ;
     RECT  1425.7 675.68 1440.86 704.44 ;
     RECT  1432.22 715.58 1440.86 723.76 ;
     RECT  1436.54 553.88 1441.34 554.08 ;
     RECT  1426.66 564.8 1441.34 565 ;
     RECT  1432.22 1022.6 1441.34 1026.58 ;
     RECT  1440.1 1183.88 1441.54 1216 ;
     RECT  1439.42 636.62 1442.02 647.74 ;
     RECT  1440.38 952.88 1442.02 953.08 ;
     RECT  1440.86 675.68 1442.3 723.76 ;
     RECT  1435.78 980.18 1442.3 980.38 ;
     RECT  1433.86 1292.24 1442.3 1300.42 ;
     RECT  1440.38 765.14 1442.5 785.08 ;
     RECT  1428.58 1131.38 1442.5 1131.58 ;
     RECT  1435.78 992.36 1442.98 992.56 ;
     RECT  1437.7 600.92 1443.46 607.42 ;
     RECT  1442.5 775.64 1443.46 785.08 ;
     RECT  1440.58 795.38 1444.42 795.58 ;
     RECT  1425.5 426.62 1444.7 426.82 ;
     RECT  1434.14 848.72 1444.7 849.34 ;
     RECT  1441.34 553.88 1444.9 565 ;
     RECT  1442.3 675.68 1444.9 724.18 ;
     RECT  1438.46 863.42 1445.18 863.62 ;
     RECT  1443.46 775.64 1445.38 775.84 ;
     RECT  1441.54 1183.88 1445.38 1212.64 ;
     RECT  1440.1 1225.46 1445.66 1227.76 ;
     RECT  1444.9 564.8 1445.86 565 ;
     RECT  1437.02 822.26 1445.86 840.1 ;
     RECT  1444.7 886.1 1446.14 886.3 ;
     RECT  1445.86 822.26 1446.62 837.58 ;
     RECT  1446.14 761.36 1446.82 761.56 ;
     RECT  1441.34 1015.46 1446.82 1032.46 ;
     RECT  1414.46 480.8 1447.1 489.4 ;
     RECT  1446.62 819.32 1447.3 837.58 ;
     RECT  1427.9 1097.78 1447.3 1116.04 ;
     RECT  1443.26 618.56 1447.58 618.76 ;
     RECT  1444.9 553.88 1447.78 554.08 ;
     RECT  1444.9 715.58 1447.78 724.18 ;
     RECT  1438.66 912.14 1448.26 928.72 ;
     RECT  1442.3 973.46 1448.26 980.38 ;
     RECT  1437.7 584.12 1448.54 592.3 ;
     RECT  1443.46 600.92 1448.54 605.74 ;
     RECT  1448.54 584.12 1448.74 605.74 ;
     RECT  1444.9 675.68 1448.74 704.44 ;
     RECT  1447.3 826.04 1448.74 837.58 ;
     RECT  1447.58 618.56 1449.02 624.64 ;
     RECT  1445.38 1183.88 1449.22 1184.08 ;
     RECT  1411.3 448.04 1449.5 448.24 ;
     RECT  1439.62 526.16 1449.5 531.82 ;
     RECT  1448.74 591.68 1449.7 605.74 ;
     RECT  1449.02 618.56 1449.7 625.06 ;
     RECT  1449.02 805.88 1449.7 806.08 ;
     RECT  1448.74 829.4 1449.7 837.58 ;
     RECT  1444.7 426.62 1449.98 433.12 ;
     RECT  1449.5 443.84 1450.18 448.24 ;
     RECT  1449.7 618.56 1450.18 618.76 ;
     RECT  1449.7 837.38 1450.18 837.58 ;
     RECT  1444.7 848.72 1450.18 853.54 ;
     RECT  1448.54 952.04 1450.18 952.24 ;
     RECT  1445.18 863.42 1450.46 864.46 ;
     RECT  1448.54 875.6 1450.46 875.8 ;
     RECT  1448.54 961.7 1450.46 961.9 ;
     RECT  1447.78 715.58 1450.66 717.04 ;
     RECT  1450.46 863.42 1450.66 875.8 ;
     RECT  1450.46 796.64 1451.14 796.84 ;
     RECT  1450.18 848.72 1451.14 849.76 ;
     RECT  1450.66 863.42 1451.14 867.4 ;
     RECT  1445.38 1196.06 1451.14 1212.64 ;
     RECT  1451.14 867.2 1451.62 867.4 ;
     RECT  1446.82 1017.56 1451.62 1032.46 ;
     RECT  1448.26 980.18 1451.9 980.38 ;
     RECT  1451.14 849.14 1452.1 849.76 ;
     RECT  1446.14 886.1 1452.1 890.08 ;
     RECT  1442.02 636.62 1452.38 640.18 ;
     RECT  1447.58 998.66 1452.58 998.86 ;
     RECT  1451.42 509.36 1453.54 509.56 ;
     RECT  1452.1 886.1 1453.54 886.3 ;
     RECT  1451.62 1017.98 1453.54 1032.46 ;
     RECT  1451.9 980.18 1454.02 984.58 ;
     RECT  1453.54 1017.98 1454.5 1026.58 ;
     RECT  1451.9 1045.28 1454.5 1045.48 ;
     RECT  1440.1 1240.58 1454.5 1271.02 ;
     RECT  1445.66 1223.78 1454.78 1227.76 ;
     RECT  1454.5 1240.58 1454.78 1244.98 ;
     RECT  1444.22 1139.36 1455.46 1139.56 ;
     RECT  1454.78 1223.78 1455.46 1244.98 ;
     RECT  1448.26 919.28 1455.94 928.72 ;
     RECT  1448.74 675.68 1456.42 692.68 ;
     RECT  1447.58 939.86 1456.42 940.06 ;
     RECT  1450.46 954.14 1456.42 961.9 ;
     RECT  1447.3 1097.78 1456.9 1108.48 ;
     RECT  1443.46 784.88 1457.38 785.08 ;
     RECT  1448.74 704.24 1457.86 704.44 ;
     RECT  1432.7 1150.7 1457.86 1150.9 ;
     RECT  1456.42 675.68 1458.34 686.8 ;
     RECT  1442.3 1290.56 1458.34 1300.42 ;
     RECT  1430.3 465.68 1458.62 470.92 ;
     RECT  1458.34 682.82 1458.82 686.8 ;
     RECT  1456.42 954.14 1459.78 954.34 ;
     RECT  1454.02 984.38 1459.78 984.58 ;
     RECT  1451.14 1196.06 1459.78 1211.8 ;
     RECT  1458.62 459.38 1460.26 470.92 ;
     RECT  1448.06 1309.88 1460.26 1310.08 ;
     RECT  1450.66 715.58 1461.22 715.78 ;
     RECT  1455.94 924.32 1461.22 928.72 ;
     RECT  1456.9 1105.76 1461.22 1108.48 ;
     RECT  1455.74 1120.46 1461.22 1120.66 ;
     RECT  1459.78 1196.06 1461.5 1199.2 ;
     RECT  1449.98 426.62 1461.7 433.54 ;
     RECT  1455.46 1223.78 1461.7 1227.76 ;
     RECT  1455.46 1240.58 1461.7 1244.98 ;
     RECT  1447.1 480.8 1462.66 497.38 ;
     RECT  1454.5 1022.6 1462.94 1026.58 ;
     RECT  1457.18 1036.46 1462.94 1036.66 ;
     RECT  1459.58 999.5 1464.1 999.7 ;
     RECT  1463.9 722.3 1464.38 722.5 ;
     RECT  1449.5 519.44 1464.58 531.82 ;
     RECT  1461.7 432.92 1465.34 433.54 ;
     RECT  1460.26 465.68 1465.34 470.92 ;
     RECT  1449.7 591.68 1465.34 602.8 ;
     RECT  1462.66 489.2 1465.54 497.38 ;
     RECT  1464.58 519.44 1465.82 519.64 ;
     RECT  1450.18 443.84 1466.78 444.04 ;
     RECT  1462.94 1022.6 1466.78 1036.66 ;
     RECT  1466.3 1045.28 1466.78 1045.48 ;
     RECT  1458.34 1294.76 1467.74 1300.42 ;
     RECT  1466.78 443.84 1468.9 444.46 ;
     RECT  1461.5 1190.18 1469.18 1199.2 ;
     RECT  1461.5 666.86 1469.66 667.06 ;
     RECT  1468.22 979.76 1469.66 979.96 ;
     RECT  1466.78 1022.6 1470.62 1045.48 ;
     RECT  1464.58 531.62 1470.82 531.82 ;
     RECT  1452.38 636.62 1470.82 640.6 ;
     RECT  1469.66 979.76 1470.82 980.38 ;
     RECT  1454.5 1256.54 1470.82 1271.02 ;
     RECT  1470.62 1015.04 1471.1 1045.48 ;
     RECT  1471.1 1010.84 1472.06 1045.48 ;
     RECT  1470.82 979.76 1472.74 979.96 ;
     RECT  1465.34 465.68 1473.02 471.34 ;
     RECT  1458.82 682.82 1473.7 683.02 ;
     RECT  1472.06 1010.84 1473.7 1045.9 ;
     RECT  1465.34 591.68 1473.98 610.78 ;
     RECT  1461.22 1105.76 1474.46 1105.96 ;
     RECT  1470.62 569 1475.14 569.2 ;
     RECT  1474.94 685.76 1475.42 685.96 ;
     RECT  1440.1 1173.8 1475.42 1174 ;
     RECT  1469.18 1188.92 1475.42 1199.2 ;
     RECT  1473.98 591.68 1475.62 617.92 ;
     RECT  1469.66 666.44 1475.9 667.06 ;
     RECT  1464.38 722.3 1475.9 728.8 ;
     RECT  1474.46 1105.76 1476.1 1109.74 ;
     RECT  1475.9 666.44 1477.34 670.42 ;
     RECT  1475.42 1173.8 1477.54 1199.2 ;
     RECT  1461.7 1241.42 1477.82 1244.98 ;
     RECT  1477.34 666.44 1478.02 671.68 ;
     RECT  1475.9 719.78 1478.5 728.8 ;
     RECT  1476.86 537.08 1478.98 537.28 ;
     RECT  1478.02 666.44 1478.98 669.58 ;
     RECT  1461.22 928.52 1479.74 928.72 ;
     RECT  1464.38 417.8 1480.9 418 ;
     RECT  1468.9 444.26 1480.9 444.46 ;
     RECT  1473.02 465.68 1481.38 475.12 ;
     RECT  1463.42 553.04 1481.86 553.24 ;
     RECT  1465.54 489.2 1482.14 489.4 ;
     RECT  1465.34 432.92 1482.82 434.38 ;
     RECT  1479.74 928.52 1482.82 932.08 ;
     RECT  1478.98 666.44 1483.3 667.06 ;
     RECT  1470.82 636.62 1483.58 640.18 ;
     RECT  1472.06 704.66 1484.74 704.86 ;
     RECT  1471.58 1309.88 1484.74 1310.08 ;
     RECT  1475.42 685.76 1486.66 691.84 ;
     RECT  1483.58 636.62 1486.94 641.02 ;
     RECT  1482.82 928.52 1487.42 928.72 ;
     RECT  1459.78 1211.6 1487.62 1211.8 ;
     RECT  1483.3 666.44 1489.06 666.64 ;
     RECT  1482.82 432.92 1489.82 433.54 ;
     RECT  1477.54 1190.18 1489.82 1199.2 ;
     RECT  1465.82 519.02 1490.3 519.64 ;
     RECT  1489.34 939.44 1490.3 939.64 ;
     RECT  1482.14 489.2 1490.5 497.38 ;
     RECT  1481.38 466.52 1490.78 475.12 ;
     RECT  1486.94 636.62 1491.26 643.96 ;
     RECT  1473.7 1010.84 1491.46 1026.58 ;
     RECT  1490.78 530.78 1491.94 530.98 ;
     RECT  1491.26 636.62 1492.42 644.38 ;
     RECT  1491.46 1010.84 1492.42 1014.82 ;
     RECT  1490.3 512.3 1492.7 519.64 ;
     RECT  1487.42 928.1 1493.66 928.72 ;
     RECT  1490.3 939.44 1493.66 943 ;
     RECT  1473.7 1037.72 1494.34 1045.9 ;
     RECT  1477.54 1173.8 1494.62 1174 ;
     RECT  1489.82 1184.72 1494.62 1199.2 ;
     RECT  1492.7 512.3 1494.82 527.62 ;
     RECT  1494.62 1173.8 1494.82 1199.2 ;
     RECT  1494.34 1037.72 1495.3 1037.92 ;
     RECT  1467.74 1294.76 1496.26 1300.84 ;
     RECT  1491.26 1150.28 1496.74 1150.48 ;
     RECT  1492.42 1010.84 1497.22 1011.04 ;
     RECT  1491.26 1135.58 1498.18 1135.78 ;
     RECT  1494.82 519.44 1498.66 527.62 ;
     RECT  1475.62 591.68 1498.94 610.78 ;
     RECT  1493.18 569 1499.42 569.2 ;
     RECT  1493.66 928.1 1499.42 943 ;
     RECT  1492.42 636.62 1499.62 643.96 ;
     RECT  1499.42 926.84 1500.1 943 ;
     RECT  1489.82 428.72 1500.58 433.54 ;
     RECT  1499.42 569 1500.58 569.62 ;
     RECT  1493.66 984.8 1500.58 985 ;
     RECT  1486.66 691.64 1501.06 691.84 ;
     RECT  1477.82 1241.42 1501.06 1245.82 ;
     RECT  1500.1 942.8 1501.34 943 ;
     RECT  1494.82 1190.18 1501.34 1199.2 ;
     RECT  1498.94 590.84 1501.54 610.78 ;
     RECT  1498.66 519.44 1502.02 521.74 ;
     RECT  1501.54 591.68 1502.5 610.78 ;
     RECT  1410.82 747.92 1502.78 748.12 ;
     RECT  1490.78 458.96 1502.98 475.12 ;
     RECT  1502.5 595.04 1502.98 610.78 ;
     RECT  1494.82 1173.8 1503.46 1177.36 ;
     RECT  1502.98 595.04 1503.94 606.58 ;
     RECT  1478.5 722.3 1503.94 728.8 ;
     RECT  1503.46 1175.9 1504.42 1177.36 ;
     RECT  1504.42 1177.16 1505.86 1177.36 ;
     RECT  1501.34 1190.18 1506.14 1202.14 ;
     RECT  1505.66 530.78 1506.34 530.98 ;
     RECT  1505.66 503.9 1506.62 504.52 ;
     RECT  1505.18 621.92 1506.62 622.12 ;
     RECT  1502.98 466.52 1506.82 475.12 ;
     RECT  1506.62 621.08 1506.82 622.12 ;
     RECT  1437 -70 1507 178 ;
     RECT  1437 1622 1507 1870 ;
     RECT  1490.78 1218.74 1507.3 1218.94 ;
     RECT  1506.14 1190.18 1507.58 1203.82 ;
     RECT  1506.82 621.08 1508.26 621.28 ;
     RECT  1486.46 1159.52 1508.26 1159.72 ;
     RECT  1490.5 489.2 1508.54 489.4 ;
     RECT  1507.58 1190.18 1508.74 1204.24 ;
     RECT  1508.74 1199 1509.22 1204.24 ;
     RECT  1506.62 500.54 1510.18 504.52 ;
     RECT  1502.02 519.44 1510.18 519.64 ;
     RECT  1500.1 926.84 1511.14 928.72 ;
     RECT  1501.34 942.8 1511.14 943.42 ;
     RECT  1511.14 942.8 1511.62 943 ;
     RECT  1505.66 992.36 1511.62 992.56 ;
     RECT  1506.82 467.36 1512.1 475.12 ;
     RECT  1510.18 503.9 1512.1 504.52 ;
     RECT  1500.58 569 1512.1 569.2 ;
     RECT  1503.94 722.3 1512.1 727.54 ;
     RECT  1502.78 746.66 1512.1 748.12 ;
     RECT  1508.74 1190.18 1512.1 1190.38 ;
     RECT  1500.58 432.92 1514.3 433.54 ;
     RECT  1512.1 467.36 1515.94 467.56 ;
     RECT  1499.62 636.62 1517.66 639.76 ;
     RECT  1511.9 616.88 1518.62 617.08 ;
     RECT  1518.62 616.88 1519.1 617.5 ;
     RECT  1517.66 632.84 1519.1 639.76 ;
     RECT  1503.94 602.6 1519.58 606.58 ;
     RECT  1515.74 1166.24 1521.5 1166.44 ;
     RECT  1514.78 663.5 1523.42 663.7 ;
     RECT  1521.5 1161.62 1523.42 1166.44 ;
     RECT  1523.42 1159.52 1524.38 1166.44 ;
     RECT  1507 0 1525 178 ;
     RECT  1507 1622 1525 1800 ;
     RECT  1523.42 663.5 1525.82 670.42 ;
     RECT  1521.02 1187.66 1526.02 1187.86 ;
     RECT  1507.1 455.6 1526.5 455.8 ;
     RECT  1518.14 518.18 1526.5 518.38 ;
     RECT  1526.3 716.42 1526.78 716.62 ;
     RECT  1519.58 602.6 1528.7 607.42 ;
     RECT  1509.22 1199 1529.18 1202.14 ;
     RECT  1525.34 689.96 1530.14 690.16 ;
     RECT  1529.18 1199 1530.14 1202.56 ;
     RECT  1528.7 601.34 1530.62 607.42 ;
     RECT  1519.1 616.88 1530.62 639.76 ;
     RECT  1530.62 555.14 1532.06 555.34 ;
     RECT  1530.62 601.34 1533.02 639.76 ;
     RECT  1525.82 663.5 1533.02 675.04 ;
     RECT  1461.7 1227.56 1533.5 1227.76 ;
     RECT  1533.02 660.56 1533.98 675.04 ;
     RECT  1530.14 686.18 1533.98 690.16 ;
     RECT  1526.78 716.42 1533.98 721.24 ;
     RECT  1533.02 600.5 1534.46 639.76 ;
     RECT  1511.9 650.06 1534.46 650.26 ;
     RECT  1533.98 660.56 1534.46 690.16 ;
     RECT  1523.42 704.66 1534.46 704.86 ;
     RECT  1533.5 1227.56 1534.46 1229.02 ;
     RECT  1501.06 1241.42 1534.46 1244.98 ;
     RECT  1514.3 432.08 1535.19 433.54 ;
     RECT  1533.98 463.16 1535.19 463.36 ;
     RECT  1531.58 474.08 1535.19 474.28 ;
     RECT  1508.54 488.78 1535.19 489.4 ;
     RECT  1532.06 554.72 1535.19 557.86 ;
     RECT  1526.3 584.12 1535.19 584.32 ;
     RECT  1534.46 595.46 1535.19 639.76 ;
     RECT  1534.46 650.06 1535.19 704.86 ;
     RECT  1533.98 715.16 1535.19 721.24 ;
     RECT  1522.46 734.9 1535.19 735.1 ;
     RECT  1512.1 747.92 1535.19 748.12 ;
     RECT  1511.14 928.52 1535.19 928.72 ;
     RECT  1491.46 1026.38 1535.19 1026.58 ;
     RECT  1404.81 1061.66 1535.19 1061.86 ;
     RECT  1476.1 1105.76 1535.19 1105.96 ;
     RECT  1524.38 1159.52 1535.19 1174 ;
     RECT  1530.14 1197.74 1535.19 1202.56 ;
     RECT  1532.54 1215.8 1535.19 1216 ;
     RECT  1534.46 1227.56 1535.19 1244.98 ;
     RECT  1470.82 1259.48 1535.19 1271.02 ;
     RECT  1496.26 1294.76 1535.19 1294.96 ;
     RECT  1535.19 215.36 1540.81 1583.92 ;
     RECT  1540.81 474.08 1541.38 474.28 ;
     RECT  1540.81 554.72 1541.38 555.34 ;
     RECT  1540.81 426.2 1541.86 436.9 ;
     RECT  1540.81 503.48 1542.82 504.52 ;
     RECT  1541.38 555.14 1543.3 555.34 ;
     RECT  1540.81 734.9 1544.26 735.1 ;
     RECT  1541.86 432.08 1545.7 436.9 ;
     RECT  1540.81 601.34 1545.7 639.76 ;
     RECT  1545.7 601.34 1546.18 607.42 ;
     RECT  1545.7 432.92 1547.14 436.9 ;
     RECT  1540.81 448.88 1547.14 463.36 ;
     RECT  1540.81 686.18 1550.3 686.38 ;
     RECT  1540.81 704.66 1550.78 711.16 ;
     RECT  1540.81 1267.04 1551.46 1271.02 ;
     RECT  1547.14 454.76 1552.42 463.36 ;
     RECT  1545.7 617.3 1552.42 639.76 ;
     RECT  1547.14 432.92 1555.78 433.12 ;
     RECT  1542.82 504.32 1556.26 504.52 ;
     RECT  1540.81 584.12 1556.26 584.32 ;
     RECT  1540.81 663.5 1556.74 670.84 ;
     RECT  1550.3 686.18 1556.74 690.16 ;
     RECT  1550.78 704.66 1556.74 712.84 ;
     RECT  1546.18 607.22 1558.18 607.42 ;
     RECT  1552.42 617.3 1558.18 625.48 ;
     RECT  1556.74 689.96 1558.18 690.16 ;
     RECT  1554.62 561.86 1561.06 562.06 ;
     RECT  1552.42 454.76 1561.54 454.96 ;
     RECT  1556.74 663.5 1561.54 663.7 ;
     RECT  1556.74 712.64 1561.54 712.84 ;
     RECT  1557.5 546.32 1562.02 546.52 ;
     RECT  1558.18 617.3 1562.5 617.5 ;
     RECT  1563.26 726.92 1564.9 727.12 ;
     RECT  1540.81 650.06 1567.3 650.26 ;
     RECT  1567.58 557.66 1569.5 557.86 ;
     RECT  1540.81 1026.38 1569.7 1026.58 ;
     RECT  1569.5 557.66 1570.18 562.48 ;
     RECT  1540.81 1294.76 1573.54 1294.96 ;
     RECT  1540.81 1199 1574.5 1199.2 ;
     RECT  1552.42 636.62 1575.46 639.76 ;
     RECT  1570.18 562.28 1576.42 562.48 ;
     RECT  1540.81 1227.56 1576.9 1227.76 ;
     RECT  1551.46 1267.04 1576.9 1267.24 ;
     RECT  1540.81 1241.42 1577.38 1244.98 ;
     RECT  1577.38 1244.78 1577.86 1244.98 ;
     RECT  1575.46 636.62 1579.3 636.82 ;
     RECT  1540.81 489.2 1588.14 489.4 ;
     RECT  1540.81 747.92 1588.14 748.12 ;
     RECT  1565.66 807.98 1588.14 808.18 ;
     RECT  1540.81 928.52 1588.14 928.72 ;
     RECT  1540.81 1061.66 1588.14 1061.86 ;
     RECT  1540.81 1105.76 1588.14 1105.96 ;
     RECT  1525 -70 1595 178 ;
     RECT  1525 1622 1595 1870 ;
     RECT  1588.14 215.36 1597.86 1583.92 ;
     RECT  1595 0 1620 178 ;
     RECT  1595 1622 1620 1800 ;
     RECT  1620 0 1622 180 ;
     RECT  1597.86 219.14 1622 1580.14 ;
     RECT  1620 1620 1622 1800 ;
     RECT  1622 0 1800 1800 ;
     RECT  1800 205 1870 275 ;
     RECT  1800 293 1870 363 ;
     RECT  1800 381 1870 451 ;
     RECT  1800 469 1870 539 ;
     RECT  1800 557 1870 627 ;
     RECT  1800 645 1870 715 ;
     RECT  1800 733 1870 803 ;
     RECT  1800 821 1870 891 ;
     RECT  1800 909 1870 979 ;
     RECT  1800 997 1870 1067 ;
     RECT  1800 1085 1870 1155 ;
     RECT  1800 1173 1870 1243 ;
     RECT  1800 1261 1870 1331 ;
     RECT  1800 1349 1870 1419 ;
     RECT  1800 1437 1870 1507 ;
     RECT  1800 1525 1870 1595 ;
    LAYER Metal5 ;
     RECT  205 -70 275 0 ;
     RECT  293 -70 363 0 ;
     RECT  381 -70 451 0 ;
     RECT  469 -70 539 0 ;
     RECT  557 -70 627 0 ;
     RECT  645 -70 715 0 ;
     RECT  733 -70 803 0 ;
     RECT  821 -70 891 0 ;
     RECT  909 -70 979 0 ;
     RECT  997 -70 1067 0 ;
     RECT  1085 -70 1155 0 ;
     RECT  1173 -70 1243 0 ;
     RECT  1261 -70 1331 0 ;
     RECT  1349 -70 1419 0 ;
     RECT  1437 -70 1507 0 ;
     RECT  1525 -70 1595 0 ;
     RECT  0 0 1800 178 ;
     RECT  0 178 180 180 ;
     RECT  1620 178 1800 180 ;
     RECT  0 180 178 205 ;
     RECT  1622 180 1800 205 ;
     RECT  1139.9 178 1140.1 215.15 ;
     RECT  -70 205 178 218.93 ;
     RECT  202.185 215.15 211.815 218.93 ;
     RECT  1185.98 178 1186.18 218.93 ;
     RECT  1406.78 178 1406.98 218.93 ;
     RECT  1588.185 215.15 1597.815 218.93 ;
     RECT  1622 205 1870 218.93 ;
     RECT  1090.46 178 1098.82 221.24 ;
     RECT  1033.82 216.2 1034.02 221.66 ;
     RECT  1018.94 220.82 1019.14 224.6 ;
     RECT  1032.86 221.66 1034.02 224.6 ;
     RECT  1054.94 178 1055.14 224.6 ;
     RECT  1068.86 197.72 1069.06 224.6 ;
     RECT  1083.26 221.24 1098.82 224.6 ;
     RECT  1185.98 218.93 1200.765 224.6 ;
     RECT  1274.3 178 1274.5 224.6 ;
     RECT  1315.58 178 1315.78 224.6 ;
     RECT  1018.94 224.6 1034.02 255.26 ;
     RECT  1052.54 224.6 1055.14 262.82 ;
     RECT  1048.22 262.82 1055.14 269.96 ;
     RECT  1068.86 224.6 1106.98 269.96 ;
     RECT  -70 218.93 211.815 275 ;
     RECT  1588.185 218.93 1870 275 ;
     RECT  0 275 211.815 293 ;
     RECT  1588.185 275 1800 293 ;
     RECT  1018.94 255.26 1037.38 334.64 ;
     RECT  1048.22 269.96 1106.98 334.64 ;
     RECT  -70 293 211.815 363 ;
     RECT  1588.185 293 1870 363 ;
     RECT  0 363 211.815 381 ;
     RECT  1588.185 363 1800 381 ;
     RECT  364.22 381.26 364.42 382.94 ;
     RECT  991.235 218.93 996.765 383.36 ;
     RECT  311.235 215.15 316.765 386.3 ;
     RECT  330.14 385.88 330.34 386.3 ;
     RECT  923.235 215.15 928.765 386.72 ;
     RECT  917.66 386.72 928.765 387.14 ;
     RECT  989.66 383.36 996.765 387.98 ;
     RECT  860.06 385.04 860.26 388.82 ;
     RECT  787.235 218.93 792.765 390.08 ;
     RECT  435.26 390.5 435.46 390.92 ;
     RECT  414.14 391.34 414.34 392.18 ;
     RECT  838.94 384.2 839.14 392.6 ;
     RECT  1018.94 334.64 1106.98 392.6 ;
     RECT  837.5 392.6 839.14 393.02 ;
     RECT  379.235 218.93 384.765 393.44 ;
     RECT  583.235 218.93 588.765 393.44 ;
     RECT  860.06 388.82 866.02 393.44 ;
     RECT  583.235 393.44 594.82 393.72 ;
     RECT  860.06 393.44 867.94 393.86 ;
     RECT  583.235 393.72 593.86 394.48 ;
     RECT  781.34 390.08 792.765 394.7 ;
     RECT  917.66 387.14 933.22 394.7 ;
     RECT  358.46 382.94 364.42 395.12 ;
     RECT  492.86 395.96 493.06 396.38 ;
     RECT  758.78 389.66 758.98 397.22 ;
     RECT  465.02 397.64 465.22 398.06 ;
     RECT  686.3 380.84 686.5 398.48 ;
     RECT  685.82 398.48 686.5 398.9 ;
     RECT  702.62 395.54 702.82 399.74 ;
     RECT  374.78 393.44 384.765 400.16 ;
     RECT  515.235 215.15 520.765 400.16 ;
     RECT  583.235 394.48 591.94 400.16 ;
     RECT  374.78 400.16 387.94 400.56 ;
     RECT  580.22 400.16 591.94 400.56 ;
     RECT  781.34 394.7 796.42 400.56 ;
     RECT  510.14 400.16 520.765 400.58 ;
     RECT  810.14 391.76 810.34 401 ;
     RECT  685.82 398.9 687.94 401.42 ;
     RECT  890.3 394.28 890.5 401.84 ;
     RECT  542.3 400.58 542.5 402.26 ;
     RECT  538.46 402.26 542.5 402.68 ;
     RECT  910.94 394.7 933.22 402.68 ;
     RECT  429.98 390.92 435.46 403.52 ;
     RECT  910.94 402.68 935.14 404.78 ;
     RECT  702.62 399.74 708.58 405.2 ;
     RECT  719.235 215.15 724.765 405.2 ;
     RECT  508.7 400.58 520.765 406.88 ;
     RECT  702.62 405.2 731.62 408.14 ;
     RECT  374.78 400.56 384.765 410.66 ;
     RECT  803.9 401 810.34 411.5 ;
     RECT  702.62 408.14 732.58 412.34 ;
     RECT  648.38 388.4 648.58 413.6 ;
     RECT  658.46 409.82 658.66 413.6 ;
     RECT  612.38 413.6 612.58 414.44 ;
     RECT  758.78 397.22 759.94 414.44 ;
     RECT  536.54 402.68 542.5 414.86 ;
     RECT  486.14 396.38 493.06 415.7 ;
     RECT  583.235 400.56 590.5 416.11 ;
     RECT  781.34 400.56 792.765 416.11 ;
     RECT  980.06 387.98 996.765 416.11 ;
     RECT  559.1 401.84 559.3 416.12 ;
     RECT  960.38 409.82 960.58 416.12 ;
     RECT  504.86 406.88 520.765 417.38 ;
     RECT  907.58 404.78 935.14 417.38 ;
     RECT  588.86 416.11 590.5 417.5 ;
     RECT  702.62 412.34 736.42 417.5 ;
     RECT  749.66 414.44 759.94 417.5 ;
     RECT  957.98 416.12 969.7 417.5 ;
     RECT  1270.46 224.6 1274.5 417.5 ;
     RECT  602.78 414.44 612.58 417.8 ;
     RECT  803.9 411.5 810.82 417.8 ;
     RECT  459.74 398.06 465.22 419.06 ;
     RECT  588.86 417.5 590.98 419.06 ;
     RECT  602.78 417.8 623.14 419.06 ;
     RECT  648.38 413.6 658.66 419.06 ;
     RECT  749.66 417.5 764.74 419.06 ;
     RECT  781.34 416.11 789.22 419.06 ;
     RECT  311.235 386.3 330.34 419.48 ;
     RECT  408.38 392.18 414.34 419.48 ;
     RECT  588.86 419.06 623.14 419.48 ;
     RECT  311.235 419.48 335.14 419.89 ;
     RECT  702.62 417.5 736.9 419.89 ;
     RECT  907.58 417.38 940.42 419.89 ;
     RECT  458.78 419.06 465.22 419.9 ;
     RECT  536.54 414.86 543.94 419.9 ;
     RECT  638.3 414.86 638.5 419.9 ;
     RECT  283.58 387.56 283.78 420.32 ;
     RECT  311.235 419.89 312.58 420.32 ;
     RECT  374.78 410.66 386.98 420.32 ;
     RECT  429.98 403.52 442.18 420.32 ;
     RECT  457.82 419.9 465.22 420.32 ;
     RECT  486.14 415.7 493.54 420.32 ;
     RECT  727.1 419.89 736.9 420.32 ;
     RECT  828.38 393.02 839.14 420.32 ;
     RECT  850.94 393.86 867.94 420.32 ;
     RECT  1013.66 392.6 1106.98 420.74 ;
     RECT  283.58 420.32 285.22 421.16 ;
     RECT  310.46 420.32 312.58 421.16 ;
     RECT  324.38 419.89 335.14 421.16 ;
     RECT  403.58 419.48 414.34 421.16 ;
     RECT  426.14 420.32 442.66 421.16 ;
     RECT  454.46 420.32 465.22 421.16 ;
     RECT  636.86 419.9 638.5 421.16 ;
     RECT  648.38 419.06 659.62 421.16 ;
     RECT  702.62 419.89 710.5 421.16 ;
     RECT  882.62 401.84 890.5 421.16 ;
     RECT  929.18 419.89 940.42 421.16 ;
     RECT  262.94 419.9 263.14 421.58 ;
     RECT  283.58 421.16 285.7 421.58 ;
     RECT  357.98 395.12 364.42 421.58 ;
     RECT  504.86 417.38 521.38 421.58 ;
     RECT  559.1 416.12 567.46 421.58 ;
     RECT  727.1 420.32 738.82 425.64 ;
     RECT  588.86 419.48 626.5 427.72 ;
     RECT  636.86 421.16 659.62 427.72 ;
     RECT  957.5 417.5 969.7 431.9 ;
     RECT  980.06 416.11 991.3 431.9 ;
     RECT  957.5 431.9 991.3 432.28 ;
     RECT  252.38 421.58 263.14 439.1 ;
     RECT  302.78 421.16 312.58 439.1 ;
     RECT  454.46 421.16 465.7 439.1 ;
     RECT  907.58 419.89 918.34 439.1 ;
     RECT  -70 381 211.815 445.555 ;
     RECT  229.34 421.58 235.3 445.555 ;
     RECT  251.9 439.1 263.14 445.555 ;
     RECT  273.5 421.58 285.7 445.555 ;
     RECT  302.3 439.1 313.06 445.555 ;
     RECT  324.38 421.16 336.1 445.555 ;
     RECT  353.18 421.58 364.42 445.555 ;
     RECT  374.3 420.32 386.98 445.555 ;
     RECT  403.58 421.16 414.82 445.555 ;
     RECT  426.14 421.16 443.14 445.555 ;
     RECT  453.98 439.1 465.7 445.555 ;
     RECT  482.3 420.32 493.54 445.555 ;
     RECT  504.38 421.58 521.38 445.555 ;
     RECT  536.54 419.9 544.42 445.555 ;
     RECT  554.78 421.58 567.46 445.555 ;
     RECT  588.86 427.72 659.62 445.555 ;
     RECT  676.7 401.42 687.94 445.555 ;
     RECT  698.78 421.16 710.5 445.555 ;
     RECT  727.1 425.64 738.34 445.555 ;
     RECT  749.18 419.06 764.74 445.555 ;
     RECT  777.5 419.06 789.22 445.555 ;
     RECT  803.9 417.8 811.78 445.555 ;
     RECT  827.9 420.32 839.62 445.555 ;
     RECT  850.46 420.32 867.94 445.555 ;
     RECT  878.78 421.16 890.5 445.555 ;
     RECT  907.1 439.1 918.34 445.555 ;
     RECT  929.18 421.16 940.9 445.555 ;
     RECT  956.54 432.28 991.3 445.555 ;
     RECT  1013.18 420.74 1106.98 445.555 ;
     RECT  -70 445.555 575.445 451 ;
     RECT  1588.185 381 1870 451 ;
     RECT  0 451 575.445 451.125 ;
     RECT  588.86 445.555 1106.98 451.125 ;
     RECT  1399.235 218.93 1406.98 453.08 ;
     RECT  229.34 451.125 575.445 456.955 ;
     RECT  588.86 451.125 994.535 456.955 ;
     RECT  0 451.125 217.46 462.525 ;
     RECT  229.34 456.955 994.535 462.525 ;
     RECT  1007.1 451.125 1106.98 462.525 ;
     RECT  1535.235 215.15 1540.765 463.16 ;
     RECT  1397.18 453.08 1406.98 465.68 ;
     RECT  0 462.525 211.815 469 ;
     RECT  1588.185 451 1800 469 ;
     RECT  956.54 462.525 991.3 471.24 ;
     RECT  1535.235 463.16 1542.82 471.76 ;
     RECT  1397.18 465.68 1412.74 480.8 ;
     RECT  749.18 462.525 764.74 489.48 ;
     RECT  403.58 462.525 414.82 489.5 ;
     RECT  957.5 471.24 991.3 489.7 ;
     RECT  1331.235 215.15 1336.765 497.18 ;
     RECT  504.38 462.525 521.38 503.16 ;
     RECT  749.18 489.48 763.3 503.16 ;
     RECT  907.1 462.525 918.34 503.9 ;
     RECT  929.18 462.525 940.9 503.9 ;
     RECT  1331.235 497.18 1337.38 503.9 ;
     RECT  504.38 503.16 517.54 504.1 ;
     RECT  907.1 503.9 940.9 512.08 ;
     RECT  -70 469 211.815 513.955 ;
     RECT  229.34 462.525 235.3 513.955 ;
     RECT  251.9 462.525 263.14 513.955 ;
     RECT  273.5 462.525 285.7 513.955 ;
     RECT  302.3 462.525 313.06 513.955 ;
     RECT  324.38 462.525 336.1 513.955 ;
     RECT  353.18 462.525 364.42 513.955 ;
     RECT  374.3 462.525 386.98 513.955 ;
     RECT  403.1 489.5 414.82 513.955 ;
     RECT  426.14 462.525 443.14 513.955 ;
     RECT  453.98 462.525 465.7 513.955 ;
     RECT  482.3 462.525 493.54 513.955 ;
     RECT  504.38 504.1 515.62 513.955 ;
     RECT  536.54 462.525 544.42 513.955 ;
     RECT  554.78 462.525 566.98 513.955 ;
     RECT  588.86 462.525 659.62 513.955 ;
     RECT  676.7 462.525 687.94 513.955 ;
     RECT  698.78 462.525 710.5 513.955 ;
     RECT  727.1 462.525 738.34 513.955 ;
     RECT  749.18 503.16 760.9 513.955 ;
     RECT  777.5 462.525 789.22 513.955 ;
     RECT  803.9 462.525 811.78 513.955 ;
     RECT  827.9 462.525 839.62 513.955 ;
     RECT  850.46 462.525 867.94 513.955 ;
     RECT  878.78 462.525 890.5 513.955 ;
     RECT  906.62 512.08 940.9 513.955 ;
     RECT  957.5 489.7 970.18 513.955 ;
     RECT  980.06 489.7 991.3 513.955 ;
     RECT  1013.18 462.525 1106.98 513.955 ;
     RECT  588.86 513.955 1106.98 518.3 ;
     RECT  -70 513.955 575.445 519.525 ;
     RECT  588.38 518.3 1106.98 519.525 ;
     RECT  229.34 519.525 575.445 525.355 ;
     RECT  588.38 519.525 994.535 525.355 ;
     RECT  1331.235 503.9 1339.3 526.58 ;
     RECT  1328.06 526.58 1339.3 527 ;
     RECT  -70 519.525 217.46 530.925 ;
     RECT  229.34 525.355 994.535 530.925 ;
     RECT  1007.1 519.525 1106.98 530.925 ;
     RECT  1505.66 503.9 1505.86 530.98 ;
     RECT  1127.235 215.15 1140.1 531.2 ;
     RECT  -70 530.925 211.815 539 ;
     RECT  1588.185 469 1870 539 ;
     RECT  907.58 530.925 940.9 541.72 ;
     RECT  957.5 530.925 991.3 541.72 ;
     RECT  1181.66 224.6 1200.765 542.12 ;
     RECT  1397.18 480.8 1414.66 542.32 ;
     RECT  1465.34 434.18 1465.54 546.32 ;
     RECT  1123.1 531.2 1140.1 549.88 ;
     RECT  676.7 530.925 687.94 551.78 ;
     RECT  229.34 530.925 235.3 551.98 ;
     RECT  251.9 530.925 263.14 551.98 ;
     RECT  273.5 530.925 285.7 551.98 ;
     RECT  302.3 530.925 313.06 551.98 ;
     RECT  324.38 530.925 336.1 551.98 ;
     RECT  353.18 530.925 364.42 551.98 ;
     RECT  374.3 530.925 386.98 551.98 ;
     RECT  403.1 530.925 415.3 551.98 ;
     RECT  426.14 530.925 443.62 551.98 ;
     RECT  453.98 530.925 465.7 551.98 ;
     RECT  482.3 530.925 493.54 551.98 ;
     RECT  536.54 530.925 544.42 551.98 ;
     RECT  588.38 530.925 659.62 551.98 ;
     RECT  675.26 551.78 687.94 551.98 ;
     RECT  698.78 530.925 710.5 551.98 ;
     RECT  749.18 530.925 760.9 551.98 ;
     RECT  850.46 530.925 868.42 551.98 ;
     RECT  878.78 530.925 890.5 551.98 ;
     RECT  907.58 541.72 991.3 551.98 ;
     RECT  233.66 551.98 233.86 552.4 ;
     RECT  285.5 551.98 285.7 552.4 ;
     RECT  305.66 551.98 313.06 552.4 ;
     RECT  330.14 551.98 335.62 552.4 ;
     RECT  358.46 551.98 363.46 552.4 ;
     RECT  374.3 551.98 385.06 552.4 ;
     RECT  984.38 551.98 991.3 552.4 ;
     RECT  362.3 552.4 363.46 552.82 ;
     RECT  486.62 551.98 493.54 552.82 ;
     RECT  537.02 551.98 544.42 552.82 ;
     RECT  675.26 551.98 687.46 552.82 ;
     RECT  699.26 551.98 710.5 552.82 ;
     RECT  850.46 551.98 866.98 552.82 ;
     RECT  430.46 551.98 442.18 553.24 ;
     RECT  537.5 552.82 544.42 553.24 ;
     RECT  588.38 551.98 633.7 553.24 ;
     RECT  675.26 552.82 681.7 553.24 ;
     RECT  911.42 551.98 968.26 553.24 ;
     RECT  675.26 553.24 675.94 553.32 ;
     RECT  617.18 553.24 633.7 553.66 ;
     RECT  617.18 553.66 619.3 554.08 ;
     RECT  588.38 553.24 602.98 554.5 ;
     RECT  727.1 530.925 738.34 554.72 ;
     RECT  1535.235 471.76 1540.765 554.72 ;
     RECT  749.18 551.98 760.42 554.92 ;
     RECT  911.42 553.24 967.3 555.34 ;
     RECT  309.5 552.4 313.06 555.35 ;
     RECT  504.38 530.925 515.62 555.35 ;
     RECT  699.74 552.82 710.5 555.35 ;
     RECT  725.18 554.72 738.34 555.35 ;
     RECT  652.22 551.98 659.14 555.6 ;
     RECT  878.78 551.98 889.06 556.18 ;
     RECT  850.46 552.82 862.18 556.6 ;
     RECT  0 539 211.815 557 ;
     RECT  1588.185 539 1800 557 ;
     RECT  554.78 530.925 566.98 557.02 ;
     RECT  588.38 554.5 602.02 557.02 ;
     RECT  827.9 530.925 839.62 557.44 ;
     RECT  403.1 551.98 412.9 557.86 ;
     RECT  777.5 530.925 789.22 558.28 ;
     RECT  588.38 557.02 601.54 559.13 ;
     RECT  782.3 558.28 789.22 559.13 ;
     RECT  991.235 552.4 991.3 559.13 ;
     RECT  1001.18 551.78 1001.38 559.13 ;
     RECT  782.3 559.13 792.765 559.34 ;
     RECT  803.9 530.925 811.78 559.34 ;
     RECT  753.98 554.92 760.42 559.54 ;
     RECT  699.74 555.35 738.34 560.38 ;
     RECT  911.42 555.34 963.46 560.8 ;
     RECT  1013.18 530.925 1106.98 561.02 ;
     RECT  537.98 553.24 544.42 561.22 ;
     RECT  912.38 560.8 963.46 561.22 ;
     RECT  1013.18 561.02 1110.34 561.44 ;
     RECT  334.46 552.4 335.62 561.64 ;
     RECT  699.74 560.38 732.1 562.06 ;
     RECT  583.235 559.13 601.54 562.48 ;
     RECT  617.18 554.08 617.38 562.48 ;
     RECT  888.38 556.18 889.06 562.48 ;
     RECT  537.98 561.22 543.94 562.9 ;
     RECT  542.3 562.9 543.94 563.32 ;
     RECT  850.46 556.6 850.66 563.74 ;
     RECT  403.1 557.86 403.78 564.16 ;
     RECT  827.9 557.44 838.66 564.58 ;
     RECT  1174.94 542.12 1200.765 564.58 ;
     RECT  782.3 559.34 811.78 565 ;
     RECT  888.38 562.48 888.58 565.42 ;
     RECT  753.98 559.54 759.46 565.84 ;
     RECT  1013.18 561.44 1115.14 566.06 ;
     RECT  1127.235 549.88 1140.1 566.06 ;
     RECT  374.3 552.4 384.765 566.48 ;
     RECT  583.235 562.48 591.94 566.48 ;
     RECT  719.235 562.06 732.1 566.68 ;
     RECT  273.98 551.98 274.18 567 ;
     RECT  374.3 566.48 387.94 567 ;
     RECT  580.22 566.48 591.94 567 ;
     RECT  784.22 565 811.78 567 ;
     RECT  491.42 552.82 492.58 567.1 ;
     RECT  832.22 564.58 838.66 567.52 ;
     RECT  921.98 561.22 963.46 567.94 ;
     RECT  1535.235 554.72 1541.38 568.36 ;
     RECT  1328.06 527 1339.78 568.58 ;
     RECT  939.74 567.94 963.46 568.7 ;
     RECT  861.02 556.6 862.18 568.78 ;
     RECT  542.3 563.32 543.46 568.9 ;
     RECT  554.78 557.02 566.02 568.9 ;
     RECT  699.74 562.06 703.3 569.62 ;
     RECT  309.5 555.35 316.765 570.04 ;
     RECT  939.74 568.7 963.94 570.04 ;
     RECT  1397.66 542.32 1414.66 570.04 ;
     RECT  543.26 568.9 543.46 570.88 ;
     RECT  1328.06 568.58 1340.26 570.88 ;
     RECT  374.3 567 384.765 571.3 ;
     RECT  959.42 570.04 963.94 571.72 ;
     RECT  753.98 565.84 758.02 571.94 ;
     RECT  1013.18 566.06 1140.1 572.56 ;
     RECT  1177.34 564.58 1200.765 572.56 ;
     RECT  457.82 551.98 465.7 572.98 ;
     RECT  752.54 571.94 758.02 572.98 ;
     RECT  504.38 555.35 520.765 573.4 ;
     RECT  991.235 559.13 1001.38 573.82 ;
     RECT  939.74 570.04 943.78 574.24 ;
     RECT  435.74 553.24 441.7 575.08 ;
     RECT  752.54 572.98 756.58 575.92 ;
     RECT  403.58 564.16 403.78 576.76 ;
     RECT  804.38 567 811.78 577.18 ;
     RECT  719.235 566.68 731.14 577.6 ;
     RECT  1013.18 572.56 1110.34 577.6 ;
     RECT  652.22 555.6 652.42 578.02 ;
     RECT  703.1 569.62 703.3 578.86 ;
     RECT  1123.1 572.56 1140.1 579.7 ;
     RECT  1461.02 546.32 1465.54 579.92 ;
     RECT  752.54 575.92 754.18 580.12 ;
     RECT  921.98 567.94 928.765 580.96 ;
     RECT  719.235 577.6 725.38 581.38 ;
     RECT  629.18 553.66 633.7 583.28 ;
     RECT  719.235 581.38 724.765 584.54 ;
     RECT  335.42 561.64 335.62 587.26 ;
     RECT  1458.14 579.92 1465.54 587.26 ;
     RECT  629.18 583.28 640.9 587.48 ;
     RECT  717.5 584.54 724.765 587.68 ;
     RECT  626.3 587.48 640.9 588.1 ;
     RECT  513.98 573.4 520.765 590.3 ;
     RECT  960.38 571.72 963.94 591.88 ;
     RECT  701.66 588.74 701.86 593.36 ;
     RECT  626.3 588.1 637.54 593.98 ;
     RECT  701.66 593.36 706.18 594.2 ;
     RECT  1535.235 568.36 1540.765 595.46 ;
     RECT  626.3 593.98 626.5 598.18 ;
     RECT  637.34 593.98 637.54 598.18 ;
     RECT  1444.7 561.44 1444.9 600.08 ;
     RECT  701.66 594.2 706.66 601.96 ;
     RECT  753.98 580.12 754.18 603.44 ;
     RECT  648.86 603.86 649.06 604.28 ;
     RECT  701.66 601.96 706.18 604.48 ;
     RECT  1534.46 595.46 1540.765 604.7 ;
     RECT  1458.14 587.26 1463.14 606.38 ;
     RECT  701.66 604.48 701.86 607 ;
     RECT  1430.78 594.62 1430.98 607.64 ;
     RECT  684.86 569 685.06 610.36 ;
     RECT  923.235 580.96 928.765 614.36 ;
     RECT  1533.98 604.7 1540.765 614.36 ;
     RECT  441.5 575.08 441.7 614.56 ;
     RECT  943.58 574.24 943.78 614.98 ;
     RECT  861.98 568.78 862.18 615.2 ;
     RECT  513.5 590.3 520.765 615.82 ;
     RECT  832.7 567.52 838.66 616.46 ;
     RECT  888.38 587.06 888.58 616.88 ;
     RECT  375.26 571.3 384.765 617.08 ;
     RECT  861.98 615.2 868.42 617.3 ;
     RECT  362.3 552.82 362.5 617.5 ;
     RECT  648.86 604.28 650.5 617.92 ;
     RECT  923.235 614.36 929.86 619.3 ;
     RECT  554.78 568.9 554.98 622.96 ;
     RECT  963.74 591.88 963.94 623.18 ;
     RECT  963.74 623.18 967.78 624.02 ;
     RECT  1399.235 570.04 1414.66 624.86 ;
     RECT  1444.7 600.08 1445.38 624.86 ;
     RECT  1458.14 606.38 1468.42 624.86 ;
     RECT  991.235 573.82 996.765 625.28 ;
     RECT  -70 557 211.815 627 ;
     RECT  1588.185 557 1870 627 ;
     RECT  1396.7 624.86 1414.66 628 ;
     RECT  787.235 567 792.765 628.36 ;
     RECT  780.38 628.36 792.765 629.26 ;
     RECT  811.58 577.18 811.78 629.48 ;
     RECT  719.235 587.68 724.765 631.16 ;
     RECT  735.26 588.32 735.46 631.16 ;
     RECT  1444.7 624.86 1468.42 632.42 ;
     RECT  991.235 625.28 997.54 634.52 ;
     RECT  753.98 603.44 760.42 634.94 ;
     RECT  491.42 567.1 491.62 635.2 ;
     RECT  583.235 567 588.765 635.2 ;
     RECT  781.34 629.26 792.765 635.2 ;
     RECT  991.235 634.52 1000.42 635.2 ;
     RECT  580.22 635.2 591.94 635.56 ;
     RECT  781.34 635.2 795.94 635.56 ;
     RECT  988.22 635.2 1001.86 635.56 ;
     RECT  1371.26 511.46 1371.46 636.82 ;
     RECT  832.22 616.46 838.66 637.46 ;
     RECT  858.62 617.3 868.42 637.88 ;
     RECT  1396.7 628 1412.74 638.5 ;
     RECT  749.18 634.94 760.42 639.98 ;
     RECT  564.86 568.9 566.02 640.4 ;
     RECT  719.235 631.16 735.46 640.4 ;
     RECT  811.58 629.48 814.18 640.4 ;
     RECT  457.82 572.98 464.26 641.86 ;
     RECT  991.235 635.56 1001.86 642.08 ;
     RECT  1013.18 577.6 1106.98 642.08 ;
     RECT  559.58 640.4 566.02 643.12 ;
     RECT  309.98 570.04 316.765 644.38 ;
     RECT  1328.06 570.88 1339.78 644.38 ;
     RECT  486.62 635.2 491.62 644.8 ;
     RECT  1530.62 614.36 1540.765 644.8 ;
     RECT  0 627 211.815 645 ;
     RECT  1588.185 627 1800 645 ;
     RECT  831.26 637.46 838.66 646.28 ;
     RECT  719.235 640.4 739.3 646.7 ;
     RECT  749.18 639.98 761.38 646.7 ;
     RECT  963.74 624.02 968.74 646.7 ;
     RECT  1426.94 607.64 1430.98 647.54 ;
     RECT  1444.22 632.42 1468.42 647.54 ;
     RECT  781.34 635.56 792.765 649.22 ;
     RECT  810.62 640.4 814.18 649.22 ;
     RECT  1399.235 638.5 1412.74 649.22 ;
     RECT  1426.94 647.54 1468.42 649.22 ;
     RECT  654.14 643.76 654.34 652.16 ;
     RECT  991.235 642.08 1106.98 653 ;
     RECT  1215.26 652.58 1215.46 653.42 ;
     RECT  653.18 652.16 654.34 655.1 ;
     RECT  704.54 653.84 704.74 655.1 ;
     RECT  940.7 655.94 940.9 656.78 ;
     RECT  957.5 646.7 968.74 656.78 ;
     RECT  515.235 615.82 520.765 657.62 ;
     RECT  311.235 644.38 316.765 658 ;
     RECT  379.235 617.08 384.765 658 ;
     RECT  583.235 635.56 588.765 658 ;
     RECT  719.235 646.7 761.38 658 ;
     RECT  923.235 619.3 929.38 658 ;
     RECT  696.86 655.1 704.74 658.04 ;
     RECT  717.98 658 761.38 658.04 ;
     RECT  262.46 551.98 262.66 658.2 ;
     RECT  513.5 657.62 522.34 658.2 ;
     RECT  309.5 658 318.34 658.24 ;
     RECT  376.22 658 387.94 658.24 ;
     RECT  580.22 658 591.94 658.24 ;
     RECT  1127.235 579.7 1140.1 658.46 ;
     RECT  853.82 637.88 868.42 658.88 ;
     RECT  696.86 658.04 761.38 659.5 ;
     RECT  921.98 658 930.34 659.72 ;
     RECT  940.7 656.78 968.74 659.72 ;
     RECT  652.7 655.1 654.34 660.56 ;
     RECT  1534.46 644.8 1540.765 660.56 ;
     RECT  681.5 659.3 681.7 662.66 ;
     RECT  696.86 659.5 734.98 662.66 ;
     RECT  1256.54 489.2 1256.74 662.66 ;
     RECT  1270.46 417.5 1274.98 662.66 ;
     RECT  921.98 659.72 968.74 663.5 ;
     RECT  668.54 659.3 668.74 663.92 ;
     RECT  681.5 662.66 734.98 663.92 ;
     RECT  745.82 659.5 761.38 665.6 ;
     RECT  515.235 658.2 522.34 666.44 ;
     RECT  652.7 660.56 657.22 667.28 ;
     RECT  668.54 663.92 734.98 667.28 ;
     RECT  849.98 658.88 868.42 667.28 ;
     RECT  878.3 665.18 878.5 667.28 ;
     RECT  907.1 655.94 907.3 667.28 ;
     RECT  917.18 663.5 968.74 667.28 ;
     RECT  745.82 665.6 770.98 667.48 ;
     RECT  849.98 667.28 878.5 667.7 ;
     RECT  888.38 616.88 891.46 667.7 ;
     RECT  559.58 643.12 565.54 669.4 ;
     RECT  583.235 658.24 588.765 669.4 ;
     RECT  1533.02 660.56 1540.765 669.58 ;
     RECT  746.3 667.48 770.98 669.8 ;
     RECT  781.34 649.22 814.18 669.8 ;
     RECT  559.58 669.4 572.26 670 ;
     RECT  583.235 669.4 590.98 670 ;
     RECT  616.7 622.34 616.9 670.22 ;
     RECT  831.26 646.28 839.62 670.64 ;
     RECT  849.98 667.7 891.46 670.64 ;
     RECT  1331.235 644.38 1339.78 670.64 ;
     RECT  1480.22 546.32 1480.42 670.84 ;
     RECT  831.26 670.64 891.46 671.06 ;
     RECT  652.7 667.28 734.98 671.26 ;
     RECT  515.235 666.44 524.74 674.84 ;
     RECT  1328.54 670.64 1339.78 675.04 ;
     RECT  1331.235 675.04 1339.78 675.46 ;
     RECT  1331.235 675.46 1338.34 675.88 ;
     RECT  1399.235 649.22 1468.42 675.88 ;
     RECT  677.18 671.26 734.98 676.1 ;
     RECT  616.7 670.22 622.18 676.52 ;
     RECT  677.18 676.1 735.94 677.36 ;
     RECT  746.3 669.8 814.18 677.36 ;
     RECT  677.18 677.36 814.18 677.98 ;
     RECT  1331.235 675.88 1337.86 677.98 ;
     RECT  652.7 671.26 663.46 678.72 ;
     RECT  605.66 673.58 605.86 681.56 ;
     RECT  1535.235 669.58 1540.765 682.4 ;
     RECT  583.235 670 588.765 683.08 ;
     RECT  652.7 678.72 662.5 683.28 ;
     RECT  580.7 683.08 591.46 683.44 ;
     RECT  544.7 687.64 546.34 688.9 ;
     RECT  601.34 681.56 605.86 688.9 ;
     RECT  652.7 683.28 660.1 689.12 ;
     RECT  542.3 692.2 544.42 692.68 ;
     RECT  581.18 683.44 590.98 692.68 ;
     RECT  1256.54 662.66 1274.98 693.32 ;
     RECT  777.5 677.98 814.18 693.52 ;
     RECT  827.9 671.06 891.46 693.74 ;
     RECT  542.3 692.68 543.94 694.36 ;
     RECT  583.235 692.68 590.98 694.48 ;
     RECT  601.34 688.9 601.54 694.48 ;
     RECT  559.58 670 565.54 695 ;
     RECT  986.3 653 1106.98 695.42 ;
     RECT  515.235 674.84 525.7 696.46 ;
     RECT  677.18 677.98 761.38 696.68 ;
     RECT  777.5 693.52 811.78 696.68 ;
     RECT  907.1 667.28 968.74 696.68 ;
     RECT  542.78 694.36 543.94 696.96 ;
     RECT  542.78 696.96 542.98 698.14 ;
     RECT  983.9 695.42 1106.98 698.36 ;
     RECT  907.1 696.68 969.22 698.78 ;
     RECT  980.54 698.36 1106.98 698.78 ;
     RECT  827.9 693.74 892.42 699.2 ;
     RECT  311.235 658.24 316.765 699.61 ;
     RECT  515.235 696.46 520.765 699.61 ;
     RECT  677.18 696.68 811.78 699.61 ;
     RECT  379.235 658.24 384.765 702.98 ;
     RECT  725.18 699.61 811.78 703.18 ;
     RECT  375.26 702.98 384.765 703.39 ;
     RECT  583.235 694.48 601.54 703.39 ;
     RECT  640.22 655.94 640.42 703.6 ;
     RECT  827.9 699.2 894.82 703.6 ;
     RECT  907.1 698.78 1106.98 703.6 ;
     RECT  273.02 703.4 281.86 703.8 ;
     RECT  593.66 703.39 601.54 703.8 ;
     RECT  1399.235 675.88 1449.22 705.5 ;
     RECT  1306.46 224.6 1315.78 708.86 ;
     RECT  1256.54 693.32 1283.62 713.48 ;
     RECT  1299.74 708.86 1315.78 713.48 ;
     RECT  -70 645 211.815 715 ;
     RECT  1588.185 645 1870 715 ;
     RECT  1398.14 705.5 1449.22 716 ;
     RECT  1533.98 682.4 1540.765 716.2 ;
     RECT  1462.94 675.88 1468.42 719.14 ;
     RECT  677.18 699.61 711.46 719.9 ;
     RECT  1181.66 572.56 1200.765 720.2 ;
     RECT  1215.26 653.42 1216.9 720.2 ;
     RECT  1370.3 659.72 1370.5 720.4 ;
     RECT  1397.66 716 1449.22 720.82 ;
     RECT  907.1 703.6 941.86 724.12 ;
     RECT  0 715 211.815 725.995 ;
     RECT  233.18 703.4 233.38 725.995 ;
     RECT  255.74 703.4 255.94 725.995 ;
     RECT  273.02 703.8 273.22 725.995 ;
     RECT  334.46 703.4 334.66 725.995 ;
     RECT  375.26 703.39 375.46 725.995 ;
     RECT  442.46 702.98 442.66 725.995 ;
     RECT  457.82 641.86 458.02 725.995 ;
     RECT  486.62 644.8 486.82 725.995 ;
     RECT  559.1 695 565.54 725.995 ;
     RECT  601.34 703.8 601.54 725.995 ;
     RECT  616.7 676.52 623.14 725.995 ;
     RECT  639.26 703.6 640.42 725.995 ;
     RECT  652.22 689.12 660.1 725.995 ;
     RECT  676.7 719.9 711.46 725.995 ;
     RECT  725.18 703.18 760.9 725.995 ;
     RECT  777.5 703.18 811.78 725.995 ;
     RECT  827.9 703.6 892.42 725.995 ;
     RECT  907.1 724.12 944.74 725.995 ;
     RECT  956.54 703.6 1106.98 725.995 ;
     RECT  0 725.995 575.445 731.565 ;
     RECT  598.105 725.995 626.455 731.565 ;
     RECT  0 731.565 217.46 733 ;
     RECT  1588.185 715 1800 733 ;
     RECT  1119.26 658.46 1140.1 734.48 ;
     RECT  1256.54 713.48 1315.78 735.74 ;
     RECT  1331.235 677.98 1336.765 735.74 ;
     RECT  1233.5 716.84 1233.7 736.16 ;
     RECT  230.025 731.565 575.445 737.395 ;
     RECT  598.105 731.565 605.855 737.395 ;
     RECT  616.7 731.565 626.455 737.395 ;
     RECT  639.26 725.995 1106.98 737.395 ;
     RECT  1398.14 720.82 1449.22 738.04 ;
     RECT  1534.46 716.2 1540.765 739.3 ;
     RECT  -70 733 217.46 742.965 ;
     RECT  230.025 737.395 581.065 742.965 ;
     RECT  592.955 737.395 605.855 742.965 ;
     RECT  616.7 737.395 1106.98 742.965 ;
     RECT  1229.66 736.16 1233.7 743.72 ;
     RECT  1168.22 741.62 1168.42 747.92 ;
     RECT  1398.14 738.04 1406.98 748.54 ;
     RECT  956.06 742.965 1106.98 750.44 ;
     RECT  1119.26 734.48 1149.22 750.44 ;
     RECT  1256.54 735.74 1336.765 751.06 ;
     RECT  1159.58 747.92 1168.42 753.8 ;
     RECT  1181.66 720.2 1216.9 753.8 ;
     RECT  1331.235 751.06 1336.765 753.8 ;
     RECT  1159.58 753.8 1216.9 755.9 ;
     RECT  676.7 742.965 760.9 756.1 ;
     RECT  956.06 750.44 1149.22 758 ;
     RECT  1159.58 755.9 1217.86 758 ;
     RECT  1468.22 719.14 1468.42 758.2 ;
     RECT  1331.235 753.8 1338.82 766.4 ;
     RECT  956.06 758 1217.86 768.08 ;
     RECT  1229.66 743.72 1238.02 768.08 ;
     RECT  956.06 768.08 1238.02 768.5 ;
     RECT  1331.235 766.4 1344.58 776.48 ;
     RECT  826.46 742.965 895.3 778.84 ;
     RECT  907.1 742.965 942.82 778.84 ;
     RECT  1418.78 738.04 1449.22 780.46 ;
     RECT  1418.78 780.46 1418.98 783.4 ;
     RECT  1355.42 761.36 1355.62 784.24 ;
     RECT  956.06 768.5 1244.26 785.3 ;
     RECT  1256.54 751.06 1320.1 785.3 ;
     RECT  777.5 742.965 811.78 785.68 ;
     RECT  826.46 778.84 942.82 787.96 ;
     RECT  956.06 785.3 1320.1 787.96 ;
     RECT  -70 742.965 211.815 794.395 ;
     RECT  233.18 742.965 233.38 794.395 ;
     RECT  255.74 742.965 255.94 794.395 ;
     RECT  334.46 742.965 334.66 794.395 ;
     RECT  375.26 742.965 375.46 794.395 ;
     RECT  442.46 742.965 442.66 794.395 ;
     RECT  457.82 742.965 458.02 794.395 ;
     RECT  486.62 742.965 486.82 794.395 ;
     RECT  559.1 742.965 565.54 794.395 ;
     RECT  601.34 742.965 601.54 794.395 ;
     RECT  616.7 742.965 623.14 794.395 ;
     RECT  639.26 742.965 640.42 794.395 ;
     RECT  652.22 742.965 660.1 794.395 ;
     RECT  676.7 756.1 715.78 794.395 ;
     RECT  727.1 756.1 760.9 794.395 ;
     RECT  777.5 785.68 815.14 794.395 ;
     RECT  826.46 787.96 1320.1 794.395 ;
     RECT  639.26 794.395 1320.1 796.64 ;
     RECT  1330.46 776.48 1344.58 796.64 ;
     RECT  1433.66 780.46 1449.22 796.64 ;
     RECT  1433.66 796.64 1450.66 798.52 ;
     RECT  -70 794.395 575.445 799.965 ;
     RECT  598.105 794.395 626.455 799.965 ;
     RECT  1380.38 758 1380.58 800 ;
     RECT  -70 799.965 217.46 803 ;
     RECT  1588.185 733 1870 803 ;
     RECT  230.025 799.965 575.445 805.795 ;
     RECT  598.105 799.965 605.855 805.795 ;
     RECT  616.7 799.965 626.455 805.795 ;
     RECT  639.26 796.64 1344.58 805.795 ;
     RECT  1449.02 798.52 1450.66 806.08 ;
     RECT  0 803 217.46 811.365 ;
     RECT  230.025 805.795 581.065 811.365 ;
     RECT  592.955 805.795 605.855 811.365 ;
     RECT  616.7 805.795 1344.58 811.365 ;
     RECT  1433.66 798.52 1438.66 818.48 ;
     RECT  1449.5 806.08 1450.66 818.48 ;
     RECT  676.7 811.365 715.78 820.9 ;
     RECT  0 811.365 211.815 821 ;
     RECT  1588.185 803 1800 821 ;
     RECT  728.06 811.365 1344.58 822.36 ;
     RECT  955.1 822.36 1344.58 824.64 ;
     RECT  957.02 824.64 1344.58 829.4 ;
     RECT  334.46 811.365 334.66 833.8 ;
     RECT  559.1 811.365 565.54 833.8 ;
     RECT  676.7 820.9 713.38 834.02 ;
     RECT  728.06 822.36 942.34 834.02 ;
     RECT  676.7 834.02 942.34 834.86 ;
     RECT  957.02 829.4 1346.98 834.86 ;
     RECT  676.7 834.86 1346.98 835.06 ;
     RECT  652.22 811.365 660.1 835.28 ;
     RECT  676.7 835.06 895.78 835.28 ;
     RECT  652.22 835.28 895.78 835.48 ;
     RECT  255.74 811.365 255.94 835.9 ;
     RECT  457.82 811.365 458.02 838 ;
     RECT  375.26 811.365 375.46 838.85 ;
     RECT  442.46 811.365 442.66 839.68 ;
     RECT  652.22 835.48 687.46 840.52 ;
     RECT  698.3 835.48 895.78 840.94 ;
     RECT  616.7 811.365 623.14 841.16 ;
     RECT  375.26 838.85 384.765 842.62 ;
     RECT  611.9 841.16 623.14 843.04 ;
     RECT  617.18 843.04 623.14 843.46 ;
     RECT  1433.66 818.48 1450.66 844.52 ;
     RECT  907.1 835.06 1346.98 845.78 ;
     RECT  704.06 840.94 895.78 847.88 ;
     RECT  906.62 845.78 1346.98 847.88 ;
     RECT  704.06 847.88 1346.98 849.14 ;
     RECT  652.7 840.52 687.46 851.44 ;
     RECT  583.235 838.85 588.765 852.5 ;
     RECT  601.34 811.365 601.54 852.5 ;
     RECT  233.18 811.365 233.38 852.92 ;
     RECT  243.26 838.64 243.46 852.92 ;
     RECT  583.235 852.5 601.54 853.34 ;
     RECT  379.235 842.62 384.765 853.76 ;
     RECT  233.18 852.92 243.46 854.28 ;
     RECT  376.22 853.76 387.94 854.28 ;
     RECT  580.22 853.34 601.54 854.28 ;
     RECT  652.7 851.44 685.06 854.38 ;
     RECT  1399.235 748.54 1406.98 856.7 ;
     RECT  653.66 854.38 685.06 857.32 ;
     RECT  704.06 849.14 1353.7 857.32 ;
     RECT  582.62 854.28 590.98 859 ;
     RECT  653.66 857.32 681.22 859.42 ;
     RECT  708.86 857.32 1353.7 859.84 ;
     RECT  242.78 854.28 243.46 860.06 ;
     RECT  673.82 859.42 681.22 860.68 ;
     RECT  639.26 811.365 640.9 861.1 ;
     RECT  1433.66 844.52 1451.14 863.62 ;
     RECT  1433.66 863.62 1449.7 864.04 ;
     RECT  653.66 859.42 663.46 864.46 ;
     RECT  1434.14 864.04 1449.7 864.46 ;
     RECT  242.78 860.06 251.62 866.36 ;
     RECT  673.82 860.68 676.9 866.98 ;
     RECT  708.86 859.84 733.54 869.08 ;
     RECT  241.82 866.36 251.62 870.98 ;
     RECT  262.46 856.28 262.66 870.98 ;
     RECT  639.26 861.1 639.46 871.6 ;
     RECT  663.26 864.46 663.46 872.86 ;
     RECT  311.235 835.07 316.765 873.49 ;
     RECT  719.235 869.08 733.54 873.49 ;
     RECT  726.14 873.49 733.54 874.76 ;
     RECT  744.38 859.84 1353.7 874.76 ;
     RECT  1434.14 864.46 1447.78 875.6 ;
     RECT  379.235 854.28 384.765 877.27 ;
     RECT  1434.14 875.6 1453.06 877.9 ;
     RECT  1380.38 800 1383.46 878.12 ;
     RECT  1397.18 856.7 1406.98 878.12 ;
     RECT  441.02 876.88 441.22 879.16 ;
     RECT  486.62 811.365 486.82 879.16 ;
     RECT  559.58 833.8 565.54 879.16 ;
     RECT  708.86 869.08 709.06 880.68 ;
     RECT  389.18 881.1 389.38 881.52 ;
     RECT  515.235 835.07 520.765 881.52 ;
     RECT  389.18 881.52 390.34 881.94 ;
     RECT  515.235 881.52 526.66 881.94 ;
     RECT  601.34 854.28 601.54 881.94 ;
     RECT  389.18 881.94 391.3 882.36 ;
     RECT  582.62 859 588.765 882.36 ;
     RECT  411.26 879.84 411.46 882.78 ;
     RECT  582.62 882.36 590.5 882.78 ;
     RECT  582.62 882.78 591.46 883.2 ;
     RECT  601.34 881.94 605.38 883.2 ;
     RECT  511.58 881.94 526.66 883.62 ;
     RECT  582.62 883.2 605.38 883.62 ;
     RECT  633.5 884.04 633.7 884.46 ;
     RECT  573.02 883.62 605.38 884.88 ;
     RECT  617.18 843.46 617.38 884.88 ;
     RECT  450.62 883.62 455.62 885.3 ;
     RECT  467.9 880.26 468.1 885.3 ;
     RECT  573.02 884.88 617.38 887.4 ;
     RECT  633.5 884.46 642.82 887.4 ;
     RECT  673.82 866.98 674.02 887.4 ;
     RECT  691.58 886.14 691.78 887.4 ;
     RECT  705.5 880.68 709.06 887.4 ;
     RECT  726.14 874.76 1353.7 887.4 ;
     RECT  691.58 887.4 693.22 889.08 ;
     RECT  411.26 882.78 412.9 889.5 ;
     RECT  450.62 885.3 470.02 889.92 ;
     RECT  491.42 885.3 496.9 890.34 ;
     RECT  705.5 887.4 1353.7 890.5 ;
     RECT  -70 821 211.815 891 ;
     RECT  1588.185 821 1870 891 ;
     RECT  1380.38 878.12 1406.98 892.82 ;
     RECT  705.5 890.5 1346.98 894.28 ;
     RECT  1380.38 892.82 1411.78 894.28 ;
     RECT  1306.46 894.28 1346.98 896.8 ;
     RECT  1331.235 896.8 1346.98 897.64 ;
     RECT  450.62 889.92 475.78 898.32 ;
     RECT  489.98 890.34 496.9 898.32 ;
     RECT  688.22 889.08 693.22 905.04 ;
     RECT  705.5 894.28 1296.58 905.04 ;
     RECT  374.3 884.04 374.5 905.46 ;
     RECT  389.18 882.36 396.1 905.46 ;
     RECT  0 891 211.815 909 ;
     RECT  1588.185 891 1800 909 ;
     RECT  1380.38 894.28 1383.46 912.76 ;
     RECT  1396.7 894.28 1411.78 916.54 ;
     RECT  573.02 887.4 674.02 923.1 ;
     RECT  1380.38 912.76 1380.58 924.94 ;
     RECT  410.3 889.5 412.9 926.46 ;
     RECT  339.74 927.72 339.94 931.08 ;
     RECT  1437.02 877.9 1453.06 943 ;
     RECT  1306.46 896.8 1321.06 943.42 ;
     RECT  688.22 905.04 1296.58 945.48 ;
     RECT  450.62 898.32 496.9 945.78 ;
     RECT  511.58 883.62 549.22 945.78 ;
     RECT  559.58 945.36 559.78 946.2 ;
     RECT  572.54 923.1 674.02 946.2 ;
     RECT  1331.235 897.64 1346.5 947.2 ;
     RECT  1438.46 943 1453.06 947.2 ;
     RECT  436.22 946.62 436.42 953.34 ;
     RECT  450.62 945.78 549.22 953.34 ;
     RECT  1399.235 916.54 1411.78 954.14 ;
     RECT  766.46 945.48 1296.58 954.34 ;
     RECT  688.22 945.48 755.62 954.6 ;
     RECT  559.58 946.2 674.02 956.9 ;
     RECT  1292.06 954.34 1296.58 957.7 ;
     RECT  1331.235 947.2 1336.765 958.34 ;
     RECT  1296.38 957.7 1296.58 958.96 ;
     RECT  1398.14 954.14 1411.78 959.18 ;
     RECT  688.22 954.6 746.5 960.22 ;
     RECT  339.74 931.08 341.86 960.48 ;
     RECT  324.86 923.94 325.06 960.9 ;
     RECT  335.42 960.48 341.86 960.9 ;
     RECT  766.46 954.34 1281.7 961.06 ;
     RECT  767.42 961.06 775.3 961.9 ;
     RECT  770.3 961.9 775.3 962.32 ;
     RECT  374.3 905.46 396.1 963.84 ;
     RECT  324.86 960.9 341.86 965.52 ;
     RECT  561.02 956.9 674.02 965.52 ;
     RECT  688.22 960.22 741.22 965.52 ;
     RECT  785.66 961.06 1281.7 965.68 ;
     RECT  436.22 953.34 549.22 967.2 ;
     RECT  561.02 965.52 741.22 967.2 ;
     RECT  324.86 965.52 347.14 969.3 ;
     RECT  436.22 967.2 741.22 970.76 ;
     RECT  773.66 962.32 775.3 972.66 ;
     RECT  785.66 965.68 1274.98 972.66 ;
     RECT  561.02 970.76 741.22 973.08 ;
     RECT  754.46 971.82 754.66 973.08 ;
     RECT  1325.66 958.34 1336.765 973.66 ;
     RECT  436.22 970.76 549.22 973.92 ;
     RECT  561.02 973.08 754.66 973.92 ;
     RECT  773.66 972.66 1274.98 973.92 ;
     RECT  374.3 963.84 400.42 976.02 ;
     RECT  1397.18 959.18 1411.78 976.82 ;
     RECT  324.86 969.3 353.38 976.86 ;
     RECT  -70 909 211.815 979 ;
     RECT  1588.185 909 1870 979 ;
     RECT  364.7 976.02 400.42 979.38 ;
     RECT  410.3 926.46 417.7 979.38 ;
     RECT  429.5 973.92 549.22 980.42 ;
     RECT  1306.46 943.42 1315.78 990.04 ;
     RECT  364.7 979.38 417.7 991.14 ;
     RECT  429.5 980.42 547.78 991.14 ;
     RECT  561.02 973.92 1274.98 992.14 ;
     RECT  364.7 991.14 547.78 992.82 ;
     RECT  363.26 992.82 547.78 994.92 ;
     RECT  561.02 992.14 1256.74 994.92 ;
     RECT  1442.78 947.2 1453.06 995.3 ;
     RECT  0 979 211.815 997 ;
     RECT  1588.185 979 1800 997 ;
     RECT  286.94 986.94 287.14 999.54 ;
     RECT  286.94 999.54 290.98 1002.06 ;
     RECT  1442.78 995.3 1453.54 1015.66 ;
     RECT  316.7 976.86 353.38 1016.34 ;
     RECT  363.26 994.92 1256.74 1016.34 ;
     RECT  1449.5 1015.66 1453.54 1017.76 ;
     RECT  1452.86 1017.76 1453.54 1018.18 ;
     RECT  1396.7 976.82 1411.78 1018.6 ;
     RECT  316.7 1016.34 1256.74 1019.48 ;
     RECT  286.94 1002.06 291.94 1021.38 ;
     RECT  278.3 1021.38 291.94 1022.22 ;
     RECT  810.62 1019.48 1256.74 1023.22 ;
     RECT  810.62 1023.22 1158.82 1023.68 ;
     RECT  316.7 1019.48 798.82 1024.52 ;
     RECT  1397.66 1018.6 1411.78 1025.74 ;
     RECT  1569.5 562.28 1569.7 1026.58 ;
     RECT  1365.5 1025.54 1365.7 1029.32 ;
     RECT  815.9 1023.68 1158.82 1029.94 ;
     RECT  1398.14 1025.74 1411.78 1029.94 ;
     RECT  1453.34 1018.18 1453.54 1032.46 ;
     RECT  316.7 1024.52 789.7 1033.34 ;
     RECT  815.9 1029.94 1152.1 1037.92 ;
     RECT  241.82 870.98 262.66 1039.02 ;
     RECT  275.42 1022.22 291.94 1039.02 ;
     RECT  1169.18 1023.22 1256.74 1044.22 ;
     RECT  758.78 1033.34 784.9 1045.1 ;
     RECT  758.78 1045.1 777.7 1047.62 ;
     RECT  1399.235 1029.94 1411.78 1048.84 ;
     RECT  316.7 1033.34 748.9 1049.3 ;
     RECT  815.9 1037.92 1096.42 1052.84 ;
     RECT  1381.34 989.42 1381.54 1055.14 ;
     RECT  1175.9 1044.22 1256.74 1058.92 ;
     RECT  1175.9 1058.92 1202.02 1060.18 ;
     RECT  1365.5 1029.32 1368.1 1066.06 ;
     RECT  -70 997 211.815 1067 ;
     RECT  1588.185 997 1870 1067 ;
     RECT  1212.38 1058.92 1256.74 1068.16 ;
     RECT  316.7 1049.3 746.98 1069.88 ;
     RECT  770.78 1047.62 777.7 1070.1 ;
     RECT  1212.38 1068.16 1214.02 1071.94 ;
     RECT  1225.34 1068.16 1256.74 1071.94 ;
     RECT  1185.98 1060.18 1202.02 1075.52 ;
     RECT  1212.38 1071.94 1212.58 1075.52 ;
     RECT  1399.235 1048.84 1404.765 1075.52 ;
     RECT  770.78 1070.1 782.02 1078.08 ;
     RECT  1235.42 1071.94 1256.74 1079.08 ;
     RECT  241.82 1039.02 291.94 1082.28 ;
     RECT  1185.98 1075.52 1212.58 1082.86 ;
     RECT  758.78 1047.62 758.98 1084.8 ;
     RECT  0 1067 211.815 1085 ;
     RECT  1588.185 1067 1800 1085 ;
     RECT  770.78 1078.08 785.86 1090.26 ;
     RECT  1175.9 1060.18 1176.1 1091.06 ;
     RECT  1306.46 990.04 1306.66 1091.26 ;
     RECT  1399.235 1075.52 1406.02 1091.9 ;
     RECT  1185.98 1082.86 1210.18 1092.52 ;
     RECT  316.7 1069.88 742.18 1092.98 ;
     RECT  758.78 1084.8 759.94 1093.2 ;
     RECT  770.78 1090.26 791.14 1093.2 ;
     RECT  1365.5 1066.06 1365.7 1093.36 ;
     RECT  1107.74 1037.92 1152.1 1094.42 ;
     RECT  1239.26 1079.08 1256.74 1094.62 ;
     RECT  758.78 1093.2 796.42 1096.76 ;
     RECT  1239.74 1094.62 1256.74 1097.98 ;
     RECT  316.7 1092.98 688.9 1098.02 ;
     RECT  1397.18 1091.9 1406.02 1098.82 ;
     RECT  1397.18 1098.82 1404.765 1099.24 ;
     RECT  765.5 1096.76 796.42 1100.76 ;
     RECT  765.5 1100.76 802.66 1101.38 ;
     RECT  1107.74 1094.42 1160.74 1101.56 ;
     RECT  1172.06 1091.06 1176.1 1101.56 ;
     RECT  241.82 1082.28 295.3 1101.6 ;
     RECT  306.62 1074.72 306.82 1101.6 ;
     RECT  1239.74 1097.98 1246.66 1101.76 ;
     RECT  316.7 1098.02 633.7 1103.9 ;
     RECT  699.74 1092.98 742.18 1103.9 ;
     RECT  772.7 1101.38 802.66 1103.9 ;
     RECT  699.74 1103.9 714.82 1104.74 ;
     RECT  1107.74 1101.56 1176.1 1105.76 ;
     RECT  1185.98 1092.52 1202.02 1105.76 ;
     RECT  645.98 1098.02 688.9 1106.42 ;
     RECT  725.18 1103.9 742.18 1107.26 ;
     RECT  779.9 1103.9 802.66 1107.26 ;
     RECT  645.98 1106.42 688.42 1108.52 ;
     RECT  649.34 1108.52 688.42 1108.94 ;
     RECT  779.9 1107.26 780.1 1111.88 ;
     RECT  560.06 1103.9 633.7 1112.3 ;
     RECT  790.94 1107.26 802.66 1112.3 ;
     RECT  815.9 1052.84 1096.9 1112.48 ;
     RECT  1107.74 1105.76 1202.02 1112.48 ;
     RECT  735.26 1107.26 742.18 1112.72 ;
     RECT  802.46 1112.3 802.66 1115.24 ;
     RECT  649.34 1108.94 686.5 1116.08 ;
     RECT  725.18 1107.26 725.38 1116.08 ;
     RECT  568.7 1112.3 633.7 1116.5 ;
     RECT  1225.34 1071.94 1225.54 1116.88 ;
     RECT  790.94 1112.3 791.14 1116.92 ;
     RECT  649.34 1116.08 651.46 1117.34 ;
     RECT  700.22 1104.74 714.82 1117.56 ;
     RECT  664.22 1116.08 686.5 1118.18 ;
     RECT  1239.74 1101.76 1245.7 1121.08 ;
     RECT  697.34 1117.56 714.82 1122.38 ;
     RECT  763.58 1120.5 763.78 1122.6 ;
     RECT  1399.235 1099.24 1404.765 1122.98 ;
     RECT  700.22 1122.38 714.82 1124.06 ;
     RECT  1245.5 1121.08 1245.7 1124.44 ;
     RECT  1397.66 1122.98 1404.765 1125.28 ;
     RECT  668.54 1118.18 686.5 1125.54 ;
     RECT  735.26 1112.72 736.9 1126.38 ;
     RECT  763.58 1122.6 766.66 1126.58 ;
     RECT  766.46 1126.58 766.66 1127 ;
     RECT  241.82 1101.6 306.82 1127.22 ;
     RECT  316.7 1103.9 547.3 1127.22 ;
     RECT  1331.235 973.66 1336.765 1128.02 ;
     RECT  651.26 1117.34 651.46 1128.48 ;
     RECT  668.54 1125.54 688.9 1128.48 ;
     RECT  730.46 1126.38 743.62 1129.1 ;
     RECT  651.26 1128.48 688.9 1130.36 ;
     RECT  633.5 1116.5 633.7 1130.58 ;
     RECT  651.26 1130.36 666.34 1130.58 ;
     RECT  815.9 1112.48 1202.02 1131.58 ;
     RECT  680.06 1130.36 688.9 1131.62 ;
     RECT  700.22 1124.06 711.94 1131.62 ;
     RECT  568.7 1116.5 618.82 1131.84 ;
     RECT  1122.62 1131.58 1202.02 1132 ;
     RECT  1173.98 1132 1202.02 1132.42 ;
     RECT  683.9 1131.62 688.9 1132.68 ;
     RECT  701.18 1131.62 711.94 1134.56 ;
     RECT  566.3 1131.84 618.82 1134.78 ;
     RECT  683.9 1132.68 689.38 1135.14 ;
     RECT  704.54 1134.56 711.94 1135.2 ;
     RECT  704.54 1135.2 713.38 1136.46 ;
     RECT  730.46 1129.1 739.3 1136.46 ;
     RECT  687.26 1135.14 689.38 1136.66 ;
     RECT  566.3 1134.78 621.7 1136.88 ;
     RECT  633.5 1130.58 666.34 1136.88 ;
     RECT  687.26 1136.66 688.42 1137.42 ;
     RECT  772.22 1137.26 772.42 1137.72 ;
     RECT  566.3 1136.88 666.34 1138.76 ;
     RECT  688.22 1137.42 688.42 1138.76 ;
     RECT  1122.62 1132 1160.74 1139.14 ;
     RECT  1122.62 1139.14 1153.06 1141.24 ;
     RECT  633.5 1138.76 666.34 1141.28 ;
     RECT  704.54 1136.46 739.3 1141.28 ;
     RECT  758.78 1137.72 772.42 1141.46 ;
     RECT  786.14 1141.04 786.34 1141.46 ;
     RECT  566.3 1138.76 621.7 1141.7 ;
     RECT  704.54 1141.28 733.06 1142.12 ;
     RECT  633.5 1141.28 657.22 1142.54 ;
     RECT  724.22 1142.12 733.06 1142.54 ;
     RECT  633.5 1142.54 645.22 1142.96 ;
     RECT  704.54 1142.12 710.5 1142.96 ;
     RECT  566.3 1141.7 618.82 1143.38 ;
     RECT  758.78 1141.46 786.34 1143.38 ;
     RECT  704.54 1142.96 710.02 1143.8 ;
     RECT  640.7 1142.96 642.34 1144.22 ;
     RECT  758.78 1143.38 760.42 1144.22 ;
     RECT  566.3 1143.38 615.94 1144.64 ;
     RECT  724.22 1142.54 724.42 1144.64 ;
     RECT  657.02 1142.54 657.22 1145.06 ;
     RECT  758.78 1144.22 758.98 1145.06 ;
     RECT  642.14 1144.22 642.34 1147.16 ;
     RECT  704.54 1143.8 704.74 1147.16 ;
     RECT  1330.46 1128.02 1336.765 1150.9 ;
     RECT  1175.9 1132.42 1202.02 1154.26 ;
     RECT  -70 1085 211.815 1155 ;
     RECT  1588.185 1085 1870 1155 ;
     RECT  241.82 1127.22 547.3 1157.66 ;
     RECT  1270.46 992.14 1274.98 1159.72 ;
     RECT  1270.94 1159.72 1274.98 1161.82 ;
     RECT  1368.86 1151.12 1369.06 1163.72 ;
     RECT  566.3 1144.64 612.58 1164.38 ;
     RECT  566.3 1164.38 605.38 1164.8 ;
     RECT  1359.74 1163.72 1369.06 1165.18 ;
     RECT  241.82 1157.66 325.54 1165.64 ;
     RECT  815.9 1131.58 1112.26 1166.24 ;
     RECT  1122.62 1141.24 1152.1 1166.24 ;
     RECT  1382.78 1162.04 1382.98 1168.96 ;
     RECT  1535.235 739.3 1540.765 1169.6 ;
     RECT  590.3 1164.8 605.38 1171.94 ;
     RECT  605.18 1171.94 605.38 1172.36 ;
     RECT  1398.14 1125.28 1404.765 1172.54 ;
     RECT  0 1155 211.815 1173 ;
     RECT  1588.185 1155 1800 1173 ;
     RECT  1398.14 1172.54 1410.82 1173.58 ;
     RECT  1399.235 1173.58 1410.82 1175.26 ;
     RECT  566.3 1164.8 576.1 1175.3 ;
     RECT  815.9 1166.24 1152.1 1177.36 ;
     RECT  590.3 1171.94 590.5 1177.82 ;
     RECT  1359.74 1165.18 1365.7 1178 ;
     RECT  815.9 1177.36 1107.94 1184.5 ;
     RECT  336.86 1157.66 547.3 1185.38 ;
     RECT  566.3 1175.3 568.9 1185.8 ;
     RECT  566.3 1185.8 566.5 1186.22 ;
     RECT  241.82 1165.64 269.38 1186.64 ;
     RECT  336.86 1185.38 536.26 1187.06 ;
     RECT  1529.66 1169.6 1540.765 1187.66 ;
     RECT  1256.54 1097.98 1256.74 1188.7 ;
     RECT  1399.235 1175.26 1404.765 1189.34 ;
     RECT  517.82 1187.06 536.26 1190 ;
     RECT  518.3 1190 536.26 1192.94 ;
     RECT  523.58 1192.94 536.26 1193.78 ;
     RECT  772.22 1143.38 786.34 1195.1 ;
     RECT  796.22 1127.6 796.42 1195.1 ;
     RECT  772.22 1195.1 796.42 1195.3 ;
     RECT  336.86 1187.06 505.06 1195.46 ;
     RECT  1118.78 1177.36 1152.1 1196.68 ;
     RECT  350.78 1195.46 505.06 1196.72 ;
     RECT  350.78 1196.72 504.1 1197.14 ;
     RECT  1398.14 1189.34 1404.765 1200.26 ;
     RECT  268.7 1186.64 269.38 1201.34 ;
     RECT  816.86 1184.5 1107.94 1202.78 ;
     RECT  336.86 1195.46 340.42 1206.6 ;
     RECT  350.78 1197.14 495.94 1206.6 ;
     RECT  816.86 1202.78 1109.38 1207.4 ;
     RECT  1119.74 1196.68 1152.1 1207.4 ;
     RECT  1455.26 1204.04 1455.46 1207.4 ;
     RECT  1439.42 1108.7 1439.62 1207.6 ;
     RECT  816.86 1207.4 1152.1 1209.7 ;
     RECT  1175.9 1154.26 1200.765 1209.7 ;
     RECT  533.18 1193.78 536.26 1210.16 ;
     RECT  816.86 1209.7 1145.86 1211.38 ;
     RECT  1331.235 1150.9 1336.765 1212.44 ;
     RECT  547.1 1185.38 547.3 1212.68 ;
     RECT  1318.46 1162.46 1318.66 1213.28 ;
     RECT  533.66 1210.16 536.26 1214.78 ;
     RECT  336.86 1206.6 495.94 1215 ;
     RECT  533.66 1214.78 534.82 1215.2 ;
     RECT  285.02 1165.64 325.54 1218.14 ;
     RECT  533.66 1215.2 533.86 1219.82 ;
     RECT  1353.98 1178 1365.7 1222.72 ;
     RECT  1185.5 1209.7 1200.765 1226.08 ;
     RECT  964.7 1211.38 1145.86 1226.5 ;
     RECT  1318.46 1213.28 1321.54 1227.98 ;
     RECT  964.7 1226.5 1142.02 1229.44 ;
     RECT  1331.235 1212.44 1337.38 1229.66 ;
     RECT  1354.46 1222.72 1365.7 1231.12 ;
     RECT  1525.82 1187.66 1540.765 1235.04 ;
     RECT  1455.26 1207.4 1459.78 1235.32 ;
     RECT  336.38 1215 495.94 1235.78 ;
     RECT  1054.46 1229.44 1142.02 1237 ;
     RECT  1166.3 1234.28 1166.5 1237.64 ;
     RECT  1270.94 1161.82 1271.14 1238.68 ;
     RECT  1530.62 1235.04 1540.765 1242.46 ;
     RECT  1054.46 1237 1141.54 1242.88 ;
     RECT  -70 1173 211.815 1243 ;
     RECT  1588.185 1173 1870 1243 ;
     RECT  1190.3 1226.08 1200.765 1244.78 ;
     RECT  1354.46 1231.12 1362.34 1245.4 ;
     RECT  1391.42 1200.26 1404.765 1245.4 ;
     RECT  293.18 1218.14 325.54 1248.18 ;
     RECT  336.38 1235.78 374.98 1248.18 ;
     RECT  964.7 1229.44 1041.22 1252.12 ;
     RECT  1166.3 1237.64 1167.46 1252.96 ;
     RECT  1331.235 1229.66 1338.82 1252.96 ;
     RECT  1459.58 1235.32 1459.78 1252.96 ;
     RECT  1190.3 1244.78 1201.54 1256.74 ;
     RECT  1192.22 1256.74 1201.54 1257.16 ;
     RECT  0 1243 211.815 1261 ;
     RECT  1588.185 1243 1800 1261 ;
     RECT  1392.38 1245.4 1404.765 1261.58 ;
     RECT  1056.38 1242.88 1141.54 1262.2 ;
     RECT  1331.235 1252.96 1337.38 1263.88 ;
     RECT  1193.66 1257.16 1201.54 1264.72 ;
     RECT  1362.14 1245.4 1362.34 1265.56 ;
     RECT  1194.14 1264.72 1201.54 1267.04 ;
     RECT  1392.38 1261.58 1405.54 1268.08 ;
     RECT  293.18 1248.18 374.98 1269.8 ;
     RECT  1167.26 1252.96 1167.46 1275.02 ;
     RECT  1331.235 1263.88 1336.765 1275.44 ;
     RECT  1119.74 1262.2 1141.54 1275.86 ;
     RECT  1156.22 1273.34 1156.42 1275.86 ;
     RECT  1166.3 1275.02 1167.46 1275.86 ;
     RECT  298.94 1269.8 374.98 1276.52 ;
     RECT  1056.38 1262.2 1106.5 1278.8 ;
     RECT  1118.3 1275.86 1141.54 1278.8 ;
     RECT  1331.235 1275.44 1337.38 1279.22 ;
     RECT  1056.38 1278.8 1141.54 1279.42 ;
     RECT  1317.98 1227.98 1321.54 1279.84 ;
     RECT  1118.3 1279.42 1141.54 1280.68 ;
     RECT  816.86 1211.38 952.42 1282.92 ;
     RECT  1392.38 1268.08 1404.765 1283.2 ;
     RECT  298.94 1276.52 325.54 1285.1 ;
     RECT  384.86 1235.78 495.94 1286.6 ;
     RECT  1194.14 1267.04 1202.02 1286.78 ;
     RECT  1194.14 1286.78 1203.46 1290.34 ;
     RECT  1331.235 1279.22 1338.82 1290.34 ;
     RECT  845.66 1282.92 952.42 1290.98 ;
     RECT  964.7 1252.12 1038.82 1290.98 ;
     RECT  1056.38 1279.42 1106.5 1292.44 ;
     RECT  1096.22 1292.44 1106.5 1292.86 ;
     RECT  336.38 1276.52 374.98 1293.74 ;
     RECT  1156.22 1275.86 1167.46 1294.96 ;
     RECT  845.66 1290.98 1038.82 1296.1 ;
     RECT  846.62 1296.1 1038.82 1297.48 ;
     RECT  269.18 1201.34 269.38 1297.94 ;
     RECT  846.62 1297.48 978.34 1298.32 ;
     RECT  341.66 1293.74 374.98 1299.62 ;
     RECT  294.62 1285.1 325.54 1301.06 ;
     RECT  341.66 1299.62 373.54 1301.3 ;
     RECT  1395.26 1283.2 1404.765 1302.52 ;
     RECT  291.26 1301.06 325.54 1304.66 ;
     RECT  988.22 1297.48 1038.82 1306.72 ;
     RECT  846.62 1298.32 952.42 1309.24 ;
     RECT  1097.18 1292.86 1106.5 1310.08 ;
     RECT  1398.14 1302.52 1404.765 1310.5 ;
     RECT  1194.62 1290.34 1203.46 1312.4 ;
     RECT  1194.62 1312.4 1203.94 1314.08 ;
     RECT  846.62 1309.24 934.66 1317.64 ;
     RECT  1119.74 1280.68 1141.54 1317.64 ;
     RECT  846.62 1317.64 931.3 1318.06 ;
     RECT  1056.38 1292.44 1082.5 1318.06 ;
     RECT  1156.22 1294.96 1166.5 1321 ;
     RECT  1194.14 1314.08 1203.94 1321 ;
     RECT  1321.34 1279.84 1321.54 1321 ;
     RECT  988.7 1306.72 1038.82 1321.42 ;
     RECT  1119.74 1317.64 1132.765 1321.84 ;
     RECT  964.7 1298.32 978.34 1322.06 ;
     RECT  988.7 1321.42 1029.7 1322.06 ;
     RECT  918.14 1318.06 931.3 1325.62 ;
     RECT  341.66 1301.3 372.58 1326.92 ;
     RECT  384.86 1286.6 490.18 1327.34 ;
     RECT  945.02 1309.24 952.42 1327.72 ;
     RECT  1156.22 1321 1156.42 1328.56 ;
     RECT  -70 1261 211.815 1331 ;
     RECT  1588.185 1261 1870 1331 ;
     RECT  341.66 1326.92 341.86 1331.96 ;
     RECT  846.62 1318.06 906.82 1332.56 ;
     RECT  846.14 1332.56 906.82 1332.88 ;
     RECT  816.86 1282.92 831.46 1333.18 ;
     RECT  844.22 1332.88 906.82 1333.18 ;
     RECT  1181.66 1308.2 1181.86 1333.6 ;
     RECT  277.82 1333.82 278.02 1335.28 ;
     RECT  422.78 1327.34 490.18 1339.1 ;
     RECT  964.7 1322.06 1029.7 1339.48 ;
     RECT  1093.82 1310.3 1094.02 1340.32 ;
     RECT  757.82 1330.46 758.02 1340.96 ;
     RECT  772.22 1195.3 795.46 1340.96 ;
     RECT  1059.26 1318.06 1082.5 1341.16 ;
     RECT  952.22 1327.72 952.42 1342.42 ;
     RECT  291.26 1304.66 317.86 1343.48 ;
     RECT  291.26 1343.48 318.82 1343.9 ;
     RECT  1127.235 1321.84 1132.765 1343.9 ;
     RECT  1195.235 1321 1203.94 1347.46 ;
     RECT  1127.235 1343.9 1134.82 1347.68 ;
     RECT  1195.235 1347.46 1202.98 1348.3 ;
     RECT  0 1331 211.815 1349 ;
     RECT  1588.185 1331 1800 1349 ;
     RECT  1073.18 1341.16 1082.5 1349.14 ;
     RECT  919.1 1325.62 931.3 1349.78 ;
     RECT  918.14 1349.78 931.3 1351.04 ;
     RECT  1040.06 1348.52 1040.26 1351.88 ;
     RECT  917.66 1351.04 931.3 1355.02 ;
     RECT  964.7 1339.48 1025.86 1357.12 ;
     RECT  384.86 1327.34 411.94 1357.58 ;
     RECT  1059.26 1341.16 1059.46 1357.96 ;
     RECT  969.5 1357.12 1025.86 1358.8 ;
     RECT  978.14 1358.8 1025.86 1359.44 ;
     RECT  917.66 1355.02 929.86 1359.64 ;
     RECT  355.1 1326.92 372.58 1360.52 ;
     RECT  978.14 1359.44 1029.7 1360.9 ;
     RECT  1127.235 1347.68 1137.22 1360.9 ;
     RECT  917.66 1359.64 928.765 1363 ;
     RECT  1040.06 1351.88 1048.42 1364.06 ;
     RECT  978.62 1360.9 1029.7 1368.46 ;
     RECT  1106.3 1310.08 1106.5 1368.46 ;
     RECT  978.62 1368.46 1016.74 1373.3 ;
     RECT  918.14 1363 928.765 1373.72 ;
     RECT  918.14 1373.72 931.78 1374.12 ;
     RECT  1097.66 1373.92 1097.86 1374.34 ;
     RECT  973.82 1373.3 1016.74 1375.18 ;
     RECT  918.14 1374.12 922.18 1375.3 ;
     RECT  982.94 1375.18 991.3 1375.3 ;
     RECT  422.78 1339.1 428.26 1377.12 ;
     RECT  438.62 1339.1 490.18 1377.12 ;
     RECT  422.78 1377.12 490.18 1379.42 ;
     RECT  355.58 1360.52 372.58 1386.32 ;
     RECT  348.86 1386.32 372.58 1387.4 ;
     RECT  384.86 1357.58 410.5 1389.08 ;
     RECT  846.62 1333.18 906.82 1396.7 ;
     RECT  918.14 1375.3 921.7 1396.7 ;
     RECT  422.78 1379.42 476.26 1406.72 ;
     RECT  1004.06 1375.18 1016.74 1407.52 ;
     RECT  439.58 1406.72 476.26 1407.56 ;
     RECT  365.18 1387.4 372.58 1411.34 ;
     RECT  441.5 1407.56 476.26 1413.02 ;
     RECT  443.42 1413.02 476.26 1414.28 ;
     RECT  422.78 1406.72 429.22 1415.54 ;
     RECT  365.18 1411.34 372.1 1418.9 ;
     RECT  -70 1349 211.815 1419 ;
     RECT  1588.185 1349 1870 1419 ;
     RECT  371.9 1418.9 372.1 1421 ;
     RECT  429.02 1415.54 429.22 1422.26 ;
     RECT  1073.18 1349.14 1073.38 1425.5 ;
     RECT  1072.7 1425.5 1073.38 1425.7 ;
     RECT  384.86 1389.08 406.66 1426.46 ;
     RECT  384.86 1426.46 390.82 1428.56 ;
     RECT  451.1 1414.28 476.26 1429.82 ;
     RECT  489.98 1379.42 490.18 1431.5 ;
     RECT  460.22 1429.82 476.26 1433.18 ;
     RECT  384.86 1428.56 385.06 1436.12 ;
     RECT  0 1419 211.815 1437 ;
     RECT  1588.185 1419 1800 1437 ;
     RECT  461.66 1433.18 476.26 1439.9 ;
     RECT  1004.06 1407.52 1006.66 1440.08 ;
     RECT  1016.54 1407.52 1016.74 1440.08 ;
     RECT  1004.06 1440.08 1016.74 1440.28 ;
     RECT  475.1 1439.9 476.26 1440.74 ;
     RECT  402.14 1426.46 406.66 1441.16 ;
     RECT  402.14 1441.16 402.34 1441.58 ;
     RECT  461.66 1439.9 461.86 1441.58 ;
     RECT  475.1 1440.74 475.3 1448.3 ;
     RECT  603.26 1449.16 605.38 1449.32 ;
     RECT  757.82 1340.96 795.46 1449.52 ;
     RECT  759.26 1449.52 795.46 1449.94 ;
     RECT  602.78 1449.32 605.86 1451.64 ;
     RECT  291.26 1343.9 323.62 1459.6 ;
     RECT  759.26 1449.94 759.46 1460.44 ;
     RECT  348.86 1387.4 349.06 1460.86 ;
     RECT  772.22 1449.94 795.46 1460.86 ;
     RECT  824.54 1333.18 831.46 1465.06 ;
     RECT  -70 1437 211.815 1507 ;
     RECT  1588.185 1437 1870 1507 ;
     RECT  917.66 1396.7 921.7 1519.24 ;
     RECT  0 1507 211.815 1525 ;
     RECT  1588.185 1507 1800 1525 ;
     RECT  831.26 1465.06 831.46 1531 ;
     RECT  845.66 1396.7 906.82 1573.42 ;
     RECT  780.86 1460.86 795.46 1577.2 ;
     RECT  921.5 1519.24 921.7 1577.2 ;
     RECT  1004.06 1440.28 1013.86 1577.2 ;
     RECT  786.14 1577.2 795.46 1577.62 ;
     RECT  851.42 1573.42 906.82 1578.04 ;
     RECT  241.82 1186.64 258.82 1578.25 ;
     RECT  294.62 1459.6 323.62 1578.25 ;
     RECT  241.82 1578.25 244.42 1578.46 ;
     RECT  311.235 1578.25 323.62 1578.46 ;
     RECT  786.14 1577.62 792.765 1578.88 ;
     RECT  895.58 1578.04 906.82 1579.3 ;
     RECT  982.94 1375.3 983.14 1579.73 ;
     RECT  -70 1525 211.815 1580.35 ;
     RECT  379.235 1579.73 384.765 1580.35 ;
     RECT  583.235 1579.73 588.765 1580.35 ;
     RECT  787.235 1578.88 792.765 1580.35 ;
     RECT  897.08 1579.3 906.82 1580.35 ;
     RECT  982.94 1579.73 996.765 1580.35 ;
     RECT  1195.235 1348.3 1200.765 1580.35 ;
     RECT  1399.235 1310.5 1404.765 1580.35 ;
     RECT  1588.185 1525 1870 1580.35 ;
     RECT  1006.46 1577.2 1013.86 1580.98 ;
     RECT  901.08 1580.35 906.82 1581.4 ;
     RECT  1026.14 1574.06 1026.34 1581.82 ;
     RECT  1072.7 1425.7 1072.9 1581.82 ;
     RECT  982.94 1580.35 983.14 1582.24 ;
     RECT  258.14 1578.25 258.82 1582.66 ;
     RECT  258.62 1582.66 258.82 1583.08 ;
     RECT  851.42 1578.04 882.34 1583.08 ;
     RECT  202.185 1580.35 211.815 1584.13 ;
     RECT  311.235 1578.46 316.765 1584.13 ;
     RECT  515.235 1583.51 520.765 1584.13 ;
     RECT  719.235 1583.51 724.765 1584.13 ;
     RECT  901.08 1581.4 902.92 1584.13 ;
     RECT  923.235 1583.51 928.765 1584.13 ;
     RECT  1127.235 1360.9 1132.765 1584.13 ;
     RECT  1331.235 1290.34 1336.765 1584.13 ;
     RECT  1535.235 1242.46 1540.765 1584.13 ;
     RECT  1588.185 1580.35 1597.815 1584.13 ;
     RECT  -70 1580.35 178 1595 ;
     RECT  1622 1580.35 1870 1595 ;
     RECT  882.14 1583.08 882.34 1601.98 ;
     RECT  1040.06 1364.06 1052.74 1603.24 ;
     RECT  0 1595 178 1620 ;
     RECT  1622 1595 1800 1620 ;
     RECT  0 1620 180 1622 ;
     RECT  964.22 1407.32 964.42 1622 ;
     RECT  1013.66 1580.98 1013.86 1622 ;
     RECT  1040.06 1603.24 1040.26 1622 ;
     RECT  1052.54 1603.24 1052.74 1622 ;
     RECT  1620 1620 1800 1622 ;
     RECT  0 1622 1800 1800 ;
     RECT  205 1800 275 1870 ;
     RECT  293 1800 363 1870 ;
     RECT  381 1800 451 1870 ;
     RECT  469 1800 539 1870 ;
     RECT  557 1800 627 1870 ;
     RECT  645 1800 715 1870 ;
     RECT  733 1800 803 1870 ;
     RECT  821 1800 891 1870 ;
     RECT  909 1800 979 1870 ;
     RECT  997 1800 1067 1870 ;
     RECT  1085 1800 1155 1870 ;
     RECT  1173 1800 1243 1870 ;
     RECT  1261 1800 1331 1870 ;
     RECT  1349 1800 1419 1870 ;
     RECT  1437 1800 1507 1870 ;
     RECT  1525 1800 1595 1870 ;
    LAYER TopMetal1 ;
     RECT  -70 205 0 1595 ;
     RECT  0 0 205 1800 ;
     RECT  205 -70 211.87 1870 ;
     RECT  211.87 725.78 272.3 743.18 ;
     RECT  211.87 513.74 273.26 531.14 ;
     RECT  261.74 657.28 280.94 658.92 ;
     RECT  272.3 721.12 280.94 743.18 ;
     RECT  211.87 -70 311.09 212 ;
     RECT  211.87 445.34 311.09 462.74 ;
     RECT  273.26 513.74 311.09 567.72 ;
     RECT  280.94 657.28 311.09 743.18 ;
     RECT  211.87 794.18 311.09 855 ;
     RECT  211.87 1588 311.09 1870 ;
     RECT  311.09 -70 316.91 462.74 ;
     RECT  311.09 513.74 316.91 743.18 ;
     RECT  311.09 794.18 316.91 874.13 ;
     RECT  311.09 1582.87 316.91 1870 ;
     RECT  316.91 -70 379.09 212 ;
     RECT  316.91 399.64 379.09 462.74 ;
     RECT  316.91 513.74 379.09 567.72 ;
     RECT  316.91 657.28 379.09 743.18 ;
     RECT  316.91 794.18 379.09 855 ;
     RECT  316.91 1588 379.09 1870 ;
     RECT  379.09 -70 384.91 462.74 ;
     RECT  379.09 513.74 384.91 743.18 ;
     RECT  379.09 794.18 384.91 877.91 ;
     RECT  379.09 1579.09 384.91 1870 ;
     RECT  384.91 794.18 440.3 855 ;
     RECT  384.91 657.28 485.9 743.18 ;
     RECT  384.91 399.64 513.26 462.74 ;
     RECT  384.91 513.74 513.26 567.72 ;
     RECT  384.91 -70 515.09 212 ;
     RECT  513.26 399.64 515.09 567.72 ;
     RECT  485.9 634.48 515.09 743.18 ;
     RECT  384.91 1588 515.09 1870 ;
     RECT  515.09 -70 520.91 743.18 ;
     RECT  515.09 1582.87 520.91 1870 ;
     RECT  520.91 399.64 522.1 567.72 ;
     RECT  440.3 794.18 577.18 877.8 ;
     RECT  520.91 -70 583.09 212 ;
     RECT  522.1 399.64 583.09 462.74 ;
     RECT  522.1 513.74 583.09 567.72 ;
     RECT  520.91 634.48 583.09 743.18 ;
     RECT  520.91 1588 583.09 1870 ;
     RECT  583.09 -70 588.91 462.74 ;
     RECT  583.09 513.74 588.91 743.18 ;
     RECT  583.09 1579.09 588.91 1870 ;
     RECT  577.18 794.18 594.82 882.36 ;
     RECT  588.91 399.64 610.22 462.74 ;
     RECT  588.91 513.74 610.22 567.72 ;
     RECT  610.22 399.64 623.86 567.72 ;
     RECT  623.86 399.64 625.3 467.4 ;
     RECT  588.91 634.48 704.3 743.18 ;
     RECT  594.82 794.18 704.3 877.8 ;
     RECT  588.91 -70 719.09 212 ;
     RECT  625.3 399.64 719.09 462.74 ;
     RECT  623.86 513.74 719.09 567.72 ;
     RECT  704.3 634.48 719.09 877.8 ;
     RECT  588.91 1588 719.09 1870 ;
     RECT  719.09 -70 724.91 462.74 ;
     RECT  719.09 513.74 724.91 877.8 ;
     RECT  719.09 1582.87 724.91 1870 ;
     RECT  724.91 634.48 736.66 877.8 ;
     RECT  736.66 721.12 751.82 877.8 ;
     RECT  750.86 930.88 754.7 932.52 ;
     RECT  751.82 721.12 756.14 882.36 ;
     RECT  754.7 930.88 756.14 955.32 ;
     RECT  756.14 721.12 784.46 955.32 ;
     RECT  724.91 -70 787.09 212 ;
     RECT  724.91 399.64 787.09 462.74 ;
     RECT  724.91 513.74 787.09 567.72 ;
     RECT  736.66 634.48 787.09 658.92 ;
     RECT  784.46 716.56 787.09 955.32 ;
     RECT  724.91 1588 787.09 1870 ;
     RECT  787.09 513.74 791.66 955.32 ;
     RECT  787.09 -70 792.91 462.74 ;
     RECT  791.66 513.74 792.91 969 ;
     RECT  787.09 1579.09 792.91 1870 ;
     RECT  792.91 721.12 819.98 969 ;
     RECT  831.5 1225 839.18 1226.64 ;
     RECT  839.18 1225 846.86 1231.2 ;
     RECT  846.86 1225 847.34 1235.76 ;
     RECT  838.22 1282 847.34 1283.64 ;
     RECT  847.34 1225 858.1 1283.64 ;
     RECT  858.1 1225 858.58 1235.76 ;
     RECT  819.98 721.12 859.06 971.28 ;
     RECT  858.58 1229.56 859.06 1235.76 ;
     RECT  859.06 1229.56 860.02 1231.2 ;
     RECT  792.91 399.64 867.7 462.74 ;
     RECT  859.06 721.12 876.82 884.64 ;
     RECT  792.91 1588 897.05 1870 ;
     RECT  897.05 1579.09 901.05 1870 ;
     RECT  901.05 1371.19 902.95 1870 ;
     RECT  792.91 513.74 915.02 567.72 ;
     RECT  792.91 -70 923.09 212 ;
     RECT  867.7 445.34 923.09 462.74 ;
     RECT  915.02 509.08 923.09 567.72 ;
     RECT  792.91 634.48 923.09 658.92 ;
     RECT  876.82 721.12 923.09 880.08 ;
     RECT  859.06 962.8 923.09 971.28 ;
     RECT  858.1 1282 923.09 1283.64 ;
     RECT  902.95 1371.19 923.09 1374.84 ;
     RECT  923.09 -70 928.91 462.74 ;
     RECT  923.09 509.08 928.91 1374.84 ;
     RECT  902.95 1582.87 928.91 1870 ;
     RECT  928.91 716.56 937.3 832.2 ;
     RECT  928.91 431.56 955.82 462.74 ;
     RECT  928.91 509.08 955.82 567.72 ;
     RECT  955.82 431.56 965.14 567.72 ;
     RECT  937.3 716.56 966.1 823.08 ;
     RECT  966.1 716.56 974.26 747.84 ;
     RECT  928.91 -70 991.09 212 ;
     RECT  965.14 431.56 991.09 462.74 ;
     RECT  965.14 513.74 991.09 567.72 ;
     RECT  928.91 634.48 991.09 658.92 ;
     RECT  974.26 716.56 991.09 743.18 ;
     RECT  966.1 794.18 991.09 823.08 ;
     RECT  928.91 960.52 991.09 962.16 ;
     RECT  928.91 1373.2 991.09 1374.84 ;
     RECT  928.91 1588 991.09 1870 ;
     RECT  991.09 -70 996.91 462.74 ;
     RECT  991.09 513.74 996.91 743.18 ;
     RECT  991.09 794.18 996.91 1374.84 ;
     RECT  991.09 1579.09 996.91 1870 ;
     RECT  996.91 445.34 1008.92 462.74 ;
     RECT  996.91 513.74 1008.92 531.14 ;
     RECT  996.91 725.78 1008.92 743.18 ;
     RECT  996.91 794.18 1008.92 811.58 ;
     RECT  1008.92 445.34 1011.52 451.34 ;
     RECT  1008.92 513.74 1011.52 519.74 ;
     RECT  1008.92 725.78 1011.52 731.78 ;
     RECT  1008.92 794.18 1011.52 800.18 ;
     RECT  996.91 634.48 1058.26 658.92 ;
     RECT  1058.26 634.48 1075.54 636.12 ;
     RECT  996.91 -70 1127.09 212 ;
     RECT  996.91 1373.2 1127.09 1374.84 ;
     RECT  996.91 1588 1127.09 1870 ;
     RECT  1127.09 -70 1132.91 1870 ;
     RECT  1132.91 -70 1195.09 212 ;
     RECT  1132.91 1588 1195.09 1870 ;
     RECT  1195.09 -70 1200.91 1870 ;
     RECT  1200.91 -70 1331.09 212 ;
     RECT  1200.91 1588 1331.09 1870 ;
     RECT  1331.09 -70 1336.91 1870 ;
     RECT  1336.91 -70 1399.09 212 ;
     RECT  1336.91 1588 1399.09 1870 ;
     RECT  1399.09 -70 1404.91 1870 ;
     RECT  1404.91 -70 1535.09 212 ;
     RECT  1404.91 1588 1535.09 1870 ;
     RECT  1535.09 -70 1540.91 1870 ;
     RECT  1540.91 -70 1588.13 212 ;
     RECT  1540.91 1588 1588.13 1870 ;
     RECT  1588.13 -70 1595 1870 ;
     RECT  1595 0 1800 1800 ;
     RECT  1800 205 1870 1595 ;
    LAYER TopMetal2 ;
     RECT  205 -70 1595 0 ;
     RECT  0 0 1800 205 ;
     RECT  -70 205 1870 212 ;
     RECT  923 212 997 1368.14 ;
     RECT  -70 212 212 1588 ;
     RECT  311 212 385 1588 ;
     RECT  515 212 589 1588 ;
     RECT  719 212 793 1588 ;
     RECT  897 1368.14 997 1588 ;
     RECT  1127 212 1201 1588 ;
     RECT  1331 212 1405 1588 ;
     RECT  1535 212 1870 1588 ;
     RECT  -70 1588 1870 1595 ;
     RECT  0 1595 1800 1800 ;
     RECT  205 1800 1595 1870 ;
  END
END croc_chip
END LIBRARY
