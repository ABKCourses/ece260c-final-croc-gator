module core_wrap (clk_i,
    core_busy_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    ref_clk_i,
    rst_ni,
    test_enable_i,
    timer0_irq_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    instr_addr_o,
    instr_rdata_i,
    irqs_i);
 input clk_i;
 output core_busy_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input ref_clk_i;
 input rst_ni;
 input test_enable_i;
 input timer0_irq_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [15:0] irqs_i;

 wire net42;
 wire net381;
 wire net378;
 wire net1048;
 wire net46;
 wire \i_ibex/branch_decision ;
 wire \i_ibex/csr_access ;
 wire \i_ibex/csr_mstatus_mie ;
 wire \i_ibex/csr_mstatus_tw ;
 wire \i_ibex/csr_mtvec_init ;
 wire \i_ibex/csr_op_en ;
 wire net72;
 wire \i_ibex/csr_restore_dret_id ;
 wire \i_ibex/csr_restore_mret_id ;
 wire \i_ibex/csr_save_cause ;
 wire \i_ibex/csr_save_id ;
 wire \i_ibex/csr_save_if ;
 wire \i_ibex/ctrl_busy ;
 wire \i_ibex/debug_csr_save ;
 wire \i_ibex/debug_ebreakm ;
 wire \i_ibex/debug_ebreaku ;
 wire \i_ibex/debug_mode ;
 wire \i_ibex/debug_single_step ;
 wire \i_ibex/div_en_ex ;
 wire \i_ibex/div_sel_ex ;
 wire \i_ibex/en_wb ;
 wire \i_ibex/ex_valid ;
 wire \i_ibex/id_in_ready ;
 wire \i_ibex/if_busy ;
 wire \i_ibex/illegal_c_insn_id ;
 wire \i_ibex/illegal_csr_insn_id ;
 wire \i_ibex/illegal_insn_id ;
 wire net254;
 wire net322;
 wire \i_ibex/instr_fetch_err ;
 wire \i_ibex/instr_fetch_err_plus2 ;
 wire \i_ibex/instr_first_cycle_id ;
 wire \i_ibex/instr_id_done ;
 wire \i_ibex/instr_is_compressed_id ;
 wire \i_ibex/instr_new_id ;
 wire \i_ibex/instr_perf_count_id ;
 wire \i_ibex/instr_req_gated ;
 wire \i_ibex/instr_valid_clear ;
 wire \i_ibex/instr_valid_id ;
 wire \i_ibex/irq_pending_o ;
 wire \i_ibex/lsu_addr_incr_req ;
 wire \i_ibex/lsu_busy ;
 wire \i_ibex/lsu_load_err ;
 wire \i_ibex/lsu_req ;
 wire \i_ibex/lsu_resp_err ;
 wire \i_ibex/lsu_resp_valid ;
 wire \i_ibex/lsu_sign_ext ;
 wire \i_ibex/lsu_store_err ;
 wire \i_ibex/lsu_we ;
 wire \i_ibex/mult_en_ex ;
 wire \i_ibex/mult_sel_ex ;
 wire \i_ibex/nmi_mode ;
 wire net1050;
 wire \i_ibex/pc_set ;
 wire \i_ibex/perf_branch ;
 wire \i_ibex/perf_div_wait ;
 wire \i_ibex/perf_dside_wait ;
 wire \i_ibex/perf_instr_ret_compressed_wb ;
 wire \i_ibex/perf_instr_ret_wb ;
 wire \i_ibex/perf_iside_wait ;
 wire \i_ibex/perf_jump ;
 wire \i_ibex/perf_load ;
 wire \i_ibex/perf_store ;
 wire \i_ibex/perf_tbranch ;
 wire \i_ibex/perf_wfi_wait ;
 wire \i_ibex/rf_ren_a ;
 wire \i_ibex/rf_ren_b ;
 wire \i_ibex/rf_we_id ;
 wire \i_ibex/rf_we_lsu ;
 wire \i_ibex/rf_we_wb ;
 wire \i_ibex/trigger_match ;
 wire \i_ibex/cs_registers_i/_0000_ ;
 wire \i_ibex/cs_registers_i/_0001_ ;
 wire \i_ibex/cs_registers_i/_0002_ ;
 wire \i_ibex/cs_registers_i/_0003_ ;
 wire \i_ibex/cs_registers_i/_0004_ ;
 wire \i_ibex/cs_registers_i/_0005_ ;
 wire net1047;
 wire net1046;
 wire net1045;
 wire net1044;
 wire \i_ibex/cs_registers_i/_0010_ ;
 wire net1043;
 wire net1042;
 wire \i_ibex/cs_registers_i/_0013_ ;
 wire net1041;
 wire net1040;
 wire \i_ibex/cs_registers_i/_0016_ ;
 wire \i_ibex/cs_registers_i/_0017_ ;
 wire net1039;
 wire net1038;
 wire \i_ibex/cs_registers_i/_0020_ ;
 wire net1037;
 wire net1036;
 wire \i_ibex/cs_registers_i/_0023_ ;
 wire net1035;
 wire \i_ibex/cs_registers_i/_0025_ ;
 wire \i_ibex/cs_registers_i/_0026_ ;
 wire \i_ibex/cs_registers_i/_0027_ ;
 wire \i_ibex/cs_registers_i/_0028_ ;
 wire net1034;
 wire net1033;
 wire net1032;
 wire \i_ibex/cs_registers_i/_0032_ ;
 wire \i_ibex/cs_registers_i/_0033_ ;
 wire net1031;
 wire net1030;
 wire \i_ibex/cs_registers_i/_0036_ ;
 wire \i_ibex/cs_registers_i/_0037_ ;
 wire \i_ibex/cs_registers_i/_0038_ ;
 wire \i_ibex/cs_registers_i/_0039_ ;
 wire \i_ibex/cs_registers_i/_0040_ ;
 wire \i_ibex/cs_registers_i/_0041_ ;
 wire \i_ibex/cs_registers_i/_0042_ ;
 wire \i_ibex/cs_registers_i/_0043_ ;
 wire \i_ibex/cs_registers_i/_0044_ ;
 wire net1029;
 wire \i_ibex/cs_registers_i/_0046_ ;
 wire \i_ibex/cs_registers_i/_0047_ ;
 wire \i_ibex/cs_registers_i/_0048_ ;
 wire \i_ibex/cs_registers_i/_0049_ ;
 wire \i_ibex/cs_registers_i/_0050_ ;
 wire \i_ibex/cs_registers_i/_0051_ ;
 wire \i_ibex/cs_registers_i/_0052_ ;
 wire \i_ibex/cs_registers_i/_0053_ ;
 wire \i_ibex/cs_registers_i/_0054_ ;
 wire \i_ibex/cs_registers_i/_0055_ ;
 wire \i_ibex/cs_registers_i/_0056_ ;
 wire \i_ibex/cs_registers_i/_0057_ ;
 wire \i_ibex/cs_registers_i/_0058_ ;
 wire \i_ibex/cs_registers_i/_0059_ ;
 wire \i_ibex/cs_registers_i/_0060_ ;
 wire \i_ibex/cs_registers_i/_0061_ ;
 wire \i_ibex/cs_registers_i/_0062_ ;
 wire \i_ibex/cs_registers_i/_0063_ ;
 wire \i_ibex/cs_registers_i/_0064_ ;
 wire \i_ibex/cs_registers_i/_0065_ ;
 wire \i_ibex/cs_registers_i/_0066_ ;
 wire \i_ibex/cs_registers_i/_0067_ ;
 wire \i_ibex/cs_registers_i/_0068_ ;
 wire \i_ibex/cs_registers_i/_0069_ ;
 wire \i_ibex/cs_registers_i/_0070_ ;
 wire \i_ibex/cs_registers_i/_0071_ ;
 wire \i_ibex/cs_registers_i/_0072_ ;
 wire \i_ibex/cs_registers_i/_0073_ ;
 wire \i_ibex/cs_registers_i/_0074_ ;
 wire \i_ibex/cs_registers_i/_0075_ ;
 wire \i_ibex/cs_registers_i/_0076_ ;
 wire \i_ibex/cs_registers_i/_0077_ ;
 wire \i_ibex/cs_registers_i/_0078_ ;
 wire \i_ibex/cs_registers_i/_0079_ ;
 wire net1028;
 wire \i_ibex/cs_registers_i/_0081_ ;
 wire \i_ibex/cs_registers_i/_0082_ ;
 wire \i_ibex/cs_registers_i/_0083_ ;
 wire \i_ibex/cs_registers_i/_0084_ ;
 wire net1027;
 wire \i_ibex/cs_registers_i/_0086_ ;
 wire \i_ibex/cs_registers_i/_0087_ ;
 wire net1026;
 wire net1025;
 wire net1024;
 wire net1023;
 wire net1022;
 wire net1021;
 wire \i_ibex/cs_registers_i/_0094_ ;
 wire net1020;
 wire net1019;
 wire \i_ibex/cs_registers_i/_0097_ ;
 wire \i_ibex/cs_registers_i/_0098_ ;
 wire \i_ibex/cs_registers_i/_0099_ ;
 wire net1018;
 wire \i_ibex/cs_registers_i/_0101_ ;
 wire \i_ibex/cs_registers_i/_0102_ ;
 wire \i_ibex/cs_registers_i/_0103_ ;
 wire \i_ibex/cs_registers_i/_0104_ ;
 wire \i_ibex/cs_registers_i/_0105_ ;
 wire \i_ibex/cs_registers_i/_0106_ ;
 wire \i_ibex/cs_registers_i/_0107_ ;
 wire \i_ibex/cs_registers_i/_0108_ ;
 wire net1017;
 wire \i_ibex/cs_registers_i/_0110_ ;
 wire \i_ibex/cs_registers_i/_0111_ ;
 wire net1016;
 wire \i_ibex/cs_registers_i/_0113_ ;
 wire \i_ibex/cs_registers_i/_0114_ ;
 wire \i_ibex/cs_registers_i/_0115_ ;
 wire \i_ibex/cs_registers_i/_0116_ ;
 wire net1015;
 wire \i_ibex/cs_registers_i/_0118_ ;
 wire net1014;
 wire \i_ibex/cs_registers_i/_0120_ ;
 wire \i_ibex/cs_registers_i/_0121_ ;
 wire \i_ibex/cs_registers_i/_0122_ ;
 wire \i_ibex/cs_registers_i/_0123_ ;
 wire \i_ibex/cs_registers_i/_0124_ ;
 wire \i_ibex/cs_registers_i/_0125_ ;
 wire net1013;
 wire \i_ibex/cs_registers_i/_0127_ ;
 wire \i_ibex/cs_registers_i/_0128_ ;
 wire \i_ibex/cs_registers_i/_0129_ ;
 wire net1012;
 wire \i_ibex/cs_registers_i/_0131_ ;
 wire net1011;
 wire \i_ibex/cs_registers_i/_0133_ ;
 wire \i_ibex/cs_registers_i/_0134_ ;
 wire \i_ibex/cs_registers_i/_0135_ ;
 wire \i_ibex/cs_registers_i/_0136_ ;
 wire net1010;
 wire net1009;
 wire net1008;
 wire \i_ibex/cs_registers_i/_0140_ ;
 wire \i_ibex/cs_registers_i/_0141_ ;
 wire net1007;
 wire net1006;
 wire \i_ibex/cs_registers_i/_0144_ ;
 wire \i_ibex/cs_registers_i/_0145_ ;
 wire \i_ibex/cs_registers_i/_0146_ ;
 wire \i_ibex/cs_registers_i/_0147_ ;
 wire \i_ibex/cs_registers_i/_0148_ ;
 wire \i_ibex/cs_registers_i/_0149_ ;
 wire \i_ibex/cs_registers_i/_0150_ ;
 wire \i_ibex/cs_registers_i/_0151_ ;
 wire net1005;
 wire \i_ibex/cs_registers_i/_0153_ ;
 wire net1004;
 wire net1003;
 wire net1002;
 wire \i_ibex/cs_registers_i/_0157_ ;
 wire net1001;
 wire \i_ibex/cs_registers_i/_0159_ ;
 wire \i_ibex/cs_registers_i/_0160_ ;
 wire \i_ibex/cs_registers_i/_0161_ ;
 wire net1000;
 wire \i_ibex/cs_registers_i/_0163_ ;
 wire \i_ibex/cs_registers_i/_0164_ ;
 wire \i_ibex/cs_registers_i/_0165_ ;
 wire net999;
 wire \i_ibex/cs_registers_i/_0167_ ;
 wire net998;
 wire \i_ibex/cs_registers_i/_0169_ ;
 wire net997;
 wire net996;
 wire net995;
 wire net994;
 wire \i_ibex/cs_registers_i/_0174_ ;
 wire \i_ibex/cs_registers_i/_0175_ ;
 wire net993;
 wire net992;
 wire net991;
 wire \i_ibex/cs_registers_i/_0179_ ;
 wire \i_ibex/cs_registers_i/_0180_ ;
 wire net990;
 wire net989;
 wire net988;
 wire \i_ibex/cs_registers_i/_0184_ ;
 wire \i_ibex/cs_registers_i/_0185_ ;
 wire \i_ibex/cs_registers_i/_0186_ ;
 wire \i_ibex/cs_registers_i/_0187_ ;
 wire \i_ibex/cs_registers_i/_0188_ ;
 wire net987;
 wire net986;
 wire \i_ibex/cs_registers_i/_0191_ ;
 wire \i_ibex/cs_registers_i/_0192_ ;
 wire \i_ibex/cs_registers_i/_0193_ ;
 wire \i_ibex/cs_registers_i/_0194_ ;
 wire \i_ibex/cs_registers_i/_0195_ ;
 wire \i_ibex/cs_registers_i/_0196_ ;
 wire \i_ibex/cs_registers_i/_0197_ ;
 wire net985;
 wire net984;
 wire \i_ibex/cs_registers_i/_0200_ ;
 wire \i_ibex/cs_registers_i/_0201_ ;
 wire \i_ibex/cs_registers_i/_0202_ ;
 wire \i_ibex/cs_registers_i/_0203_ ;
 wire \i_ibex/cs_registers_i/_0204_ ;
 wire net983;
 wire \i_ibex/cs_registers_i/_0206_ ;
 wire net982;
 wire \i_ibex/cs_registers_i/_0208_ ;
 wire net981;
 wire net980;
 wire net979;
 wire net978;
 wire \i_ibex/cs_registers_i/_0213_ ;
 wire \i_ibex/cs_registers_i/_0214_ ;
 wire net977;
 wire \i_ibex/cs_registers_i/_0216_ ;
 wire net976;
 wire \i_ibex/cs_registers_i/_0218_ ;
 wire net975;
 wire \i_ibex/cs_registers_i/_0220_ ;
 wire \i_ibex/cs_registers_i/_0221_ ;
 wire \i_ibex/cs_registers_i/_0222_ ;
 wire \i_ibex/cs_registers_i/_0223_ ;
 wire \i_ibex/cs_registers_i/_0224_ ;
 wire \i_ibex/cs_registers_i/_0225_ ;
 wire net974;
 wire \i_ibex/cs_registers_i/_0227_ ;
 wire \i_ibex/cs_registers_i/_0228_ ;
 wire net973;
 wire net972;
 wire \i_ibex/cs_registers_i/_0231_ ;
 wire \i_ibex/cs_registers_i/_0232_ ;
 wire \i_ibex/cs_registers_i/_0233_ ;
 wire \i_ibex/cs_registers_i/_0234_ ;
 wire net971;
 wire net970;
 wire \i_ibex/cs_registers_i/_0237_ ;
 wire \i_ibex/cs_registers_i/_0238_ ;
 wire \i_ibex/cs_registers_i/_0239_ ;
 wire \i_ibex/cs_registers_i/_0240_ ;
 wire \i_ibex/cs_registers_i/_0241_ ;
 wire \i_ibex/cs_registers_i/_0242_ ;
 wire \i_ibex/cs_registers_i/_0243_ ;
 wire \i_ibex/cs_registers_i/_0244_ ;
 wire \i_ibex/cs_registers_i/_0245_ ;
 wire \i_ibex/cs_registers_i/_0246_ ;
 wire \i_ibex/cs_registers_i/_0247_ ;
 wire \i_ibex/cs_registers_i/_0248_ ;
 wire \i_ibex/cs_registers_i/_0249_ ;
 wire \i_ibex/cs_registers_i/_0250_ ;
 wire \i_ibex/cs_registers_i/_0251_ ;
 wire \i_ibex/cs_registers_i/_0252_ ;
 wire \i_ibex/cs_registers_i/_0253_ ;
 wire \i_ibex/cs_registers_i/_0254_ ;
 wire \i_ibex/cs_registers_i/_0255_ ;
 wire \i_ibex/cs_registers_i/_0256_ ;
 wire \i_ibex/cs_registers_i/_0257_ ;
 wire \i_ibex/cs_registers_i/_0258_ ;
 wire \i_ibex/cs_registers_i/_0259_ ;
 wire \i_ibex/cs_registers_i/_0260_ ;
 wire \i_ibex/cs_registers_i/_0261_ ;
 wire \i_ibex/cs_registers_i/_0262_ ;
 wire \i_ibex/cs_registers_i/_0263_ ;
 wire \i_ibex/cs_registers_i/_0264_ ;
 wire \i_ibex/cs_registers_i/_0265_ ;
 wire \i_ibex/cs_registers_i/_0266_ ;
 wire \i_ibex/cs_registers_i/_0267_ ;
 wire \i_ibex/cs_registers_i/_0268_ ;
 wire \i_ibex/cs_registers_i/_0269_ ;
 wire \i_ibex/cs_registers_i/_0270_ ;
 wire \i_ibex/cs_registers_i/_0271_ ;
 wire \i_ibex/cs_registers_i/_0272_ ;
 wire \i_ibex/cs_registers_i/_0273_ ;
 wire \i_ibex/cs_registers_i/_0274_ ;
 wire \i_ibex/cs_registers_i/_0275_ ;
 wire \i_ibex/cs_registers_i/_0276_ ;
 wire \i_ibex/cs_registers_i/_0277_ ;
 wire \i_ibex/cs_registers_i/_0278_ ;
 wire \i_ibex/cs_registers_i/_0279_ ;
 wire \i_ibex/cs_registers_i/_0280_ ;
 wire \i_ibex/cs_registers_i/_0281_ ;
 wire \i_ibex/cs_registers_i/_0282_ ;
 wire \i_ibex/cs_registers_i/_0283_ ;
 wire \i_ibex/cs_registers_i/_0284_ ;
 wire \i_ibex/cs_registers_i/_0285_ ;
 wire \i_ibex/cs_registers_i/_0286_ ;
 wire \i_ibex/cs_registers_i/_0287_ ;
 wire \i_ibex/cs_registers_i/_0288_ ;
 wire \i_ibex/cs_registers_i/_0289_ ;
 wire \i_ibex/cs_registers_i/_0290_ ;
 wire \i_ibex/cs_registers_i/_0291_ ;
 wire \i_ibex/cs_registers_i/_0292_ ;
 wire \i_ibex/cs_registers_i/_0293_ ;
 wire \i_ibex/cs_registers_i/_0294_ ;
 wire \i_ibex/cs_registers_i/_0295_ ;
 wire \i_ibex/cs_registers_i/_0296_ ;
 wire \i_ibex/cs_registers_i/_0297_ ;
 wire \i_ibex/cs_registers_i/_0298_ ;
 wire \i_ibex/cs_registers_i/_0299_ ;
 wire \i_ibex/cs_registers_i/_0300_ ;
 wire \i_ibex/cs_registers_i/_0301_ ;
 wire \i_ibex/cs_registers_i/_0302_ ;
 wire \i_ibex/cs_registers_i/_0303_ ;
 wire \i_ibex/cs_registers_i/_0304_ ;
 wire \i_ibex/cs_registers_i/_0305_ ;
 wire \i_ibex/cs_registers_i/_0306_ ;
 wire \i_ibex/cs_registers_i/_0307_ ;
 wire \i_ibex/cs_registers_i/_0308_ ;
 wire \i_ibex/cs_registers_i/_0309_ ;
 wire \i_ibex/cs_registers_i/_0310_ ;
 wire \i_ibex/cs_registers_i/_0311_ ;
 wire \i_ibex/cs_registers_i/_0312_ ;
 wire \i_ibex/cs_registers_i/_0313_ ;
 wire \i_ibex/cs_registers_i/_0314_ ;
 wire \i_ibex/cs_registers_i/_0315_ ;
 wire \i_ibex/cs_registers_i/_0316_ ;
 wire \i_ibex/cs_registers_i/_0317_ ;
 wire \i_ibex/cs_registers_i/_0318_ ;
 wire \i_ibex/cs_registers_i/_0319_ ;
 wire \i_ibex/cs_registers_i/_0320_ ;
 wire \i_ibex/cs_registers_i/_0321_ ;
 wire \i_ibex/cs_registers_i/_0322_ ;
 wire \i_ibex/cs_registers_i/_0323_ ;
 wire \i_ibex/cs_registers_i/_0324_ ;
 wire \i_ibex/cs_registers_i/_0325_ ;
 wire \i_ibex/cs_registers_i/_0326_ ;
 wire \i_ibex/cs_registers_i/_0327_ ;
 wire \i_ibex/cs_registers_i/_0328_ ;
 wire \i_ibex/cs_registers_i/_0329_ ;
 wire \i_ibex/cs_registers_i/_0330_ ;
 wire \i_ibex/cs_registers_i/_0331_ ;
 wire \i_ibex/cs_registers_i/_0332_ ;
 wire \i_ibex/cs_registers_i/_0333_ ;
 wire \i_ibex/cs_registers_i/_0334_ ;
 wire \i_ibex/cs_registers_i/_0335_ ;
 wire \i_ibex/cs_registers_i/_0336_ ;
 wire \i_ibex/cs_registers_i/_0337_ ;
 wire \i_ibex/cs_registers_i/_0338_ ;
 wire \i_ibex/cs_registers_i/_0339_ ;
 wire \i_ibex/cs_registers_i/_0340_ ;
 wire net969;
 wire \i_ibex/cs_registers_i/_0342_ ;
 wire \i_ibex/cs_registers_i/_0343_ ;
 wire \i_ibex/cs_registers_i/_0344_ ;
 wire \i_ibex/cs_registers_i/_0345_ ;
 wire \i_ibex/cs_registers_i/_0346_ ;
 wire \i_ibex/cs_registers_i/_0347_ ;
 wire \i_ibex/cs_registers_i/_0348_ ;
 wire \i_ibex/cs_registers_i/_0349_ ;
 wire \i_ibex/cs_registers_i/_0350_ ;
 wire \i_ibex/cs_registers_i/_0351_ ;
 wire \i_ibex/cs_registers_i/_0352_ ;
 wire \i_ibex/cs_registers_i/_0353_ ;
 wire \i_ibex/cs_registers_i/_0354_ ;
 wire \i_ibex/cs_registers_i/_0355_ ;
 wire \i_ibex/cs_registers_i/_0356_ ;
 wire \i_ibex/cs_registers_i/_0357_ ;
 wire \i_ibex/cs_registers_i/_0358_ ;
 wire \i_ibex/cs_registers_i/_0359_ ;
 wire \i_ibex/cs_registers_i/_0360_ ;
 wire \i_ibex/cs_registers_i/_0361_ ;
 wire \i_ibex/cs_registers_i/_0362_ ;
 wire \i_ibex/cs_registers_i/_0363_ ;
 wire \i_ibex/cs_registers_i/_0364_ ;
 wire \i_ibex/cs_registers_i/_0365_ ;
 wire \i_ibex/cs_registers_i/_0366_ ;
 wire \i_ibex/cs_registers_i/_0367_ ;
 wire \i_ibex/cs_registers_i/_0368_ ;
 wire \i_ibex/cs_registers_i/_0369_ ;
 wire \i_ibex/cs_registers_i/_0370_ ;
 wire \i_ibex/cs_registers_i/_0371_ ;
 wire \i_ibex/cs_registers_i/_0372_ ;
 wire \i_ibex/cs_registers_i/_0373_ ;
 wire \i_ibex/cs_registers_i/_0374_ ;
 wire \i_ibex/cs_registers_i/_0375_ ;
 wire \i_ibex/cs_registers_i/_0376_ ;
 wire \i_ibex/cs_registers_i/_0377_ ;
 wire \i_ibex/cs_registers_i/_0378_ ;
 wire \i_ibex/cs_registers_i/_0379_ ;
 wire \i_ibex/cs_registers_i/_0380_ ;
 wire \i_ibex/cs_registers_i/_0381_ ;
 wire \i_ibex/cs_registers_i/_0382_ ;
 wire \i_ibex/cs_registers_i/_0383_ ;
 wire \i_ibex/cs_registers_i/_0384_ ;
 wire \i_ibex/cs_registers_i/_0385_ ;
 wire \i_ibex/cs_registers_i/_0386_ ;
 wire \i_ibex/cs_registers_i/_0387_ ;
 wire \i_ibex/cs_registers_i/_0388_ ;
 wire \i_ibex/cs_registers_i/_0389_ ;
 wire \i_ibex/cs_registers_i/_0390_ ;
 wire net968;
 wire net967;
 wire net966;
 wire \i_ibex/cs_registers_i/_0394_ ;
 wire net965;
 wire \i_ibex/cs_registers_i/_0396_ ;
 wire \i_ibex/cs_registers_i/_0397_ ;
 wire \i_ibex/cs_registers_i/_0398_ ;
 wire \i_ibex/cs_registers_i/_0399_ ;
 wire \i_ibex/cs_registers_i/_0400_ ;
 wire \i_ibex/cs_registers_i/_0401_ ;
 wire \i_ibex/cs_registers_i/_0402_ ;
 wire \i_ibex/cs_registers_i/_0403_ ;
 wire \i_ibex/cs_registers_i/_0404_ ;
 wire \i_ibex/cs_registers_i/_0405_ ;
 wire \i_ibex/cs_registers_i/_0406_ ;
 wire \i_ibex/cs_registers_i/_0407_ ;
 wire \i_ibex/cs_registers_i/_0408_ ;
 wire \i_ibex/cs_registers_i/_0409_ ;
 wire \i_ibex/cs_registers_i/_0410_ ;
 wire \i_ibex/cs_registers_i/_0411_ ;
 wire \i_ibex/cs_registers_i/_0412_ ;
 wire \i_ibex/cs_registers_i/_0413_ ;
 wire \i_ibex/cs_registers_i/_0414_ ;
 wire \i_ibex/cs_registers_i/_0415_ ;
 wire \i_ibex/cs_registers_i/_0416_ ;
 wire \i_ibex/cs_registers_i/_0417_ ;
 wire \i_ibex/cs_registers_i/_0418_ ;
 wire \i_ibex/cs_registers_i/_0419_ ;
 wire \i_ibex/cs_registers_i/_0420_ ;
 wire \i_ibex/cs_registers_i/_0421_ ;
 wire \i_ibex/cs_registers_i/_0422_ ;
 wire \i_ibex/cs_registers_i/_0423_ ;
 wire \i_ibex/cs_registers_i/_0424_ ;
 wire \i_ibex/cs_registers_i/_0425_ ;
 wire \i_ibex/cs_registers_i/_0426_ ;
 wire \i_ibex/cs_registers_i/_0427_ ;
 wire \i_ibex/cs_registers_i/_0428_ ;
 wire \i_ibex/cs_registers_i/_0429_ ;
 wire \i_ibex/cs_registers_i/_0430_ ;
 wire \i_ibex/cs_registers_i/_0431_ ;
 wire \i_ibex/cs_registers_i/_0432_ ;
 wire \i_ibex/cs_registers_i/_0433_ ;
 wire \i_ibex/cs_registers_i/_0434_ ;
 wire \i_ibex/cs_registers_i/_0435_ ;
 wire \i_ibex/cs_registers_i/_0436_ ;
 wire \i_ibex/cs_registers_i/_0437_ ;
 wire \i_ibex/cs_registers_i/_0438_ ;
 wire \i_ibex/cs_registers_i/_0439_ ;
 wire \i_ibex/cs_registers_i/_0440_ ;
 wire \i_ibex/cs_registers_i/_0441_ ;
 wire \i_ibex/cs_registers_i/_0442_ ;
 wire \i_ibex/cs_registers_i/_0443_ ;
 wire \i_ibex/cs_registers_i/_0444_ ;
 wire \i_ibex/cs_registers_i/_0445_ ;
 wire \i_ibex/cs_registers_i/_0446_ ;
 wire \i_ibex/cs_registers_i/_0447_ ;
 wire \i_ibex/cs_registers_i/_0448_ ;
 wire \i_ibex/cs_registers_i/_0449_ ;
 wire \i_ibex/cs_registers_i/_0450_ ;
 wire \i_ibex/cs_registers_i/_0451_ ;
 wire \i_ibex/cs_registers_i/_0452_ ;
 wire \i_ibex/cs_registers_i/_0453_ ;
 wire \i_ibex/cs_registers_i/_0454_ ;
 wire \i_ibex/cs_registers_i/_0455_ ;
 wire \i_ibex/cs_registers_i/_0456_ ;
 wire \i_ibex/cs_registers_i/_0457_ ;
 wire \i_ibex/cs_registers_i/_0458_ ;
 wire \i_ibex/cs_registers_i/_0459_ ;
 wire \i_ibex/cs_registers_i/_0460_ ;
 wire \i_ibex/cs_registers_i/_0461_ ;
 wire \i_ibex/cs_registers_i/_0462_ ;
 wire \i_ibex/cs_registers_i/_0463_ ;
 wire \i_ibex/cs_registers_i/_0464_ ;
 wire \i_ibex/cs_registers_i/_0465_ ;
 wire \i_ibex/cs_registers_i/_0466_ ;
 wire \i_ibex/cs_registers_i/_0467_ ;
 wire \i_ibex/cs_registers_i/_0468_ ;
 wire \i_ibex/cs_registers_i/_0469_ ;
 wire \i_ibex/cs_registers_i/_0470_ ;
 wire \i_ibex/cs_registers_i/_0471_ ;
 wire net964;
 wire \i_ibex/cs_registers_i/_0473_ ;
 wire \i_ibex/cs_registers_i/_0474_ ;
 wire \i_ibex/cs_registers_i/_0475_ ;
 wire \i_ibex/cs_registers_i/_0476_ ;
 wire \i_ibex/cs_registers_i/_0477_ ;
 wire \i_ibex/cs_registers_i/_0478_ ;
 wire \i_ibex/cs_registers_i/_0479_ ;
 wire \i_ibex/cs_registers_i/_0480_ ;
 wire \i_ibex/cs_registers_i/_0481_ ;
 wire \i_ibex/cs_registers_i/_0482_ ;
 wire \i_ibex/cs_registers_i/_0483_ ;
 wire \i_ibex/cs_registers_i/_0484_ ;
 wire \i_ibex/cs_registers_i/_0485_ ;
 wire \i_ibex/cs_registers_i/_0486_ ;
 wire \i_ibex/cs_registers_i/_0487_ ;
 wire \i_ibex/cs_registers_i/_0488_ ;
 wire \i_ibex/cs_registers_i/_0489_ ;
 wire \i_ibex/cs_registers_i/_0490_ ;
 wire \i_ibex/cs_registers_i/_0491_ ;
 wire \i_ibex/cs_registers_i/_0492_ ;
 wire \i_ibex/cs_registers_i/_0493_ ;
 wire \i_ibex/cs_registers_i/_0494_ ;
 wire \i_ibex/cs_registers_i/_0495_ ;
 wire \i_ibex/cs_registers_i/_0496_ ;
 wire \i_ibex/cs_registers_i/_0497_ ;
 wire \i_ibex/cs_registers_i/_0498_ ;
 wire \i_ibex/cs_registers_i/_0499_ ;
 wire \i_ibex/cs_registers_i/_0500_ ;
 wire \i_ibex/cs_registers_i/_0501_ ;
 wire \i_ibex/cs_registers_i/_0502_ ;
 wire \i_ibex/cs_registers_i/_0503_ ;
 wire \i_ibex/cs_registers_i/_0504_ ;
 wire \i_ibex/cs_registers_i/_0505_ ;
 wire \i_ibex/cs_registers_i/_0506_ ;
 wire \i_ibex/cs_registers_i/_0507_ ;
 wire \i_ibex/cs_registers_i/_0508_ ;
 wire \i_ibex/cs_registers_i/_0509_ ;
 wire \i_ibex/cs_registers_i/_0510_ ;
 wire \i_ibex/cs_registers_i/_0511_ ;
 wire \i_ibex/cs_registers_i/_0512_ ;
 wire \i_ibex/cs_registers_i/_0513_ ;
 wire \i_ibex/cs_registers_i/_0514_ ;
 wire \i_ibex/cs_registers_i/_0515_ ;
 wire \i_ibex/cs_registers_i/_0516_ ;
 wire \i_ibex/cs_registers_i/_0517_ ;
 wire \i_ibex/cs_registers_i/_0518_ ;
 wire \i_ibex/cs_registers_i/_0519_ ;
 wire \i_ibex/cs_registers_i/_0520_ ;
 wire \i_ibex/cs_registers_i/_0521_ ;
 wire \i_ibex/cs_registers_i/_0522_ ;
 wire \i_ibex/cs_registers_i/_0523_ ;
 wire \i_ibex/cs_registers_i/_0524_ ;
 wire \i_ibex/cs_registers_i/_0525_ ;
 wire \i_ibex/cs_registers_i/_0526_ ;
 wire \i_ibex/cs_registers_i/_0527_ ;
 wire \i_ibex/cs_registers_i/_0528_ ;
 wire \i_ibex/cs_registers_i/_0529_ ;
 wire \i_ibex/cs_registers_i/_0530_ ;
 wire \i_ibex/cs_registers_i/_0531_ ;
 wire \i_ibex/cs_registers_i/_0532_ ;
 wire \i_ibex/cs_registers_i/_0533_ ;
 wire \i_ibex/cs_registers_i/_0534_ ;
 wire \i_ibex/cs_registers_i/_0535_ ;
 wire \i_ibex/cs_registers_i/_0536_ ;
 wire \i_ibex/cs_registers_i/_0537_ ;
 wire \i_ibex/cs_registers_i/_0538_ ;
 wire \i_ibex/cs_registers_i/_0539_ ;
 wire \i_ibex/cs_registers_i/_0540_ ;
 wire \i_ibex/cs_registers_i/_0541_ ;
 wire \i_ibex/cs_registers_i/_0542_ ;
 wire \i_ibex/cs_registers_i/_0543_ ;
 wire \i_ibex/cs_registers_i/_0544_ ;
 wire \i_ibex/cs_registers_i/_0545_ ;
 wire \i_ibex/cs_registers_i/_0546_ ;
 wire \i_ibex/cs_registers_i/_0547_ ;
 wire \i_ibex/cs_registers_i/_0548_ ;
 wire \i_ibex/cs_registers_i/_0549_ ;
 wire \i_ibex/cs_registers_i/_0550_ ;
 wire \i_ibex/cs_registers_i/_0551_ ;
 wire \i_ibex/cs_registers_i/_0552_ ;
 wire \i_ibex/cs_registers_i/_0553_ ;
 wire \i_ibex/cs_registers_i/_0554_ ;
 wire \i_ibex/cs_registers_i/_0555_ ;
 wire \i_ibex/cs_registers_i/_0556_ ;
 wire \i_ibex/cs_registers_i/_0557_ ;
 wire \i_ibex/cs_registers_i/_0558_ ;
 wire \i_ibex/cs_registers_i/_0559_ ;
 wire \i_ibex/cs_registers_i/_0560_ ;
 wire \i_ibex/cs_registers_i/_0561_ ;
 wire \i_ibex/cs_registers_i/_0562_ ;
 wire \i_ibex/cs_registers_i/_0563_ ;
 wire \i_ibex/cs_registers_i/_0564_ ;
 wire \i_ibex/cs_registers_i/_0565_ ;
 wire \i_ibex/cs_registers_i/_0566_ ;
 wire \i_ibex/cs_registers_i/_0567_ ;
 wire \i_ibex/cs_registers_i/_0568_ ;
 wire \i_ibex/cs_registers_i/_0569_ ;
 wire \i_ibex/cs_registers_i/_0570_ ;
 wire \i_ibex/cs_registers_i/_0571_ ;
 wire \i_ibex/cs_registers_i/_0572_ ;
 wire \i_ibex/cs_registers_i/_0573_ ;
 wire \i_ibex/cs_registers_i/_0574_ ;
 wire \i_ibex/cs_registers_i/_0575_ ;
 wire \i_ibex/cs_registers_i/_0576_ ;
 wire \i_ibex/cs_registers_i/_0577_ ;
 wire \i_ibex/cs_registers_i/_0578_ ;
 wire \i_ibex/cs_registers_i/_0579_ ;
 wire \i_ibex/cs_registers_i/_0580_ ;
 wire \i_ibex/cs_registers_i/_0581_ ;
 wire \i_ibex/cs_registers_i/_0582_ ;
 wire \i_ibex/cs_registers_i/_0583_ ;
 wire \i_ibex/cs_registers_i/_0584_ ;
 wire \i_ibex/cs_registers_i/_0585_ ;
 wire \i_ibex/cs_registers_i/_0586_ ;
 wire \i_ibex/cs_registers_i/_0587_ ;
 wire \i_ibex/cs_registers_i/_0588_ ;
 wire \i_ibex/cs_registers_i/_0589_ ;
 wire \i_ibex/cs_registers_i/_0590_ ;
 wire \i_ibex/cs_registers_i/_0591_ ;
 wire \i_ibex/cs_registers_i/_0592_ ;
 wire \i_ibex/cs_registers_i/_0593_ ;
 wire net963;
 wire \i_ibex/cs_registers_i/_0595_ ;
 wire \i_ibex/cs_registers_i/_0596_ ;
 wire \i_ibex/cs_registers_i/_0597_ ;
 wire \i_ibex/cs_registers_i/_0598_ ;
 wire \i_ibex/cs_registers_i/_0599_ ;
 wire \i_ibex/cs_registers_i/_0600_ ;
 wire \i_ibex/cs_registers_i/_0601_ ;
 wire \i_ibex/cs_registers_i/_0602_ ;
 wire \i_ibex/cs_registers_i/_0603_ ;
 wire \i_ibex/cs_registers_i/_0604_ ;
 wire \i_ibex/cs_registers_i/_0605_ ;
 wire \i_ibex/cs_registers_i/_0606_ ;
 wire \i_ibex/cs_registers_i/_0607_ ;
 wire \i_ibex/cs_registers_i/_0608_ ;
 wire \i_ibex/cs_registers_i/_0609_ ;
 wire \i_ibex/cs_registers_i/_0610_ ;
 wire \i_ibex/cs_registers_i/_0611_ ;
 wire \i_ibex/cs_registers_i/_0612_ ;
 wire \i_ibex/cs_registers_i/_0613_ ;
 wire \i_ibex/cs_registers_i/_0614_ ;
 wire \i_ibex/cs_registers_i/_0615_ ;
 wire \i_ibex/cs_registers_i/_0616_ ;
 wire \i_ibex/cs_registers_i/_0617_ ;
 wire \i_ibex/cs_registers_i/_0618_ ;
 wire \i_ibex/cs_registers_i/_0619_ ;
 wire \i_ibex/cs_registers_i/_0620_ ;
 wire \i_ibex/cs_registers_i/_0621_ ;
 wire \i_ibex/cs_registers_i/_0622_ ;
 wire \i_ibex/cs_registers_i/_0623_ ;
 wire \i_ibex/cs_registers_i/_0624_ ;
 wire \i_ibex/cs_registers_i/_0625_ ;
 wire \i_ibex/cs_registers_i/_0626_ ;
 wire \i_ibex/cs_registers_i/_0627_ ;
 wire \i_ibex/cs_registers_i/_0628_ ;
 wire \i_ibex/cs_registers_i/_0629_ ;
 wire \i_ibex/cs_registers_i/_0630_ ;
 wire \i_ibex/cs_registers_i/_0631_ ;
 wire \i_ibex/cs_registers_i/_0632_ ;
 wire \i_ibex/cs_registers_i/_0633_ ;
 wire \i_ibex/cs_registers_i/_0634_ ;
 wire \i_ibex/cs_registers_i/_0635_ ;
 wire \i_ibex/cs_registers_i/_0636_ ;
 wire \i_ibex/cs_registers_i/_0637_ ;
 wire \i_ibex/cs_registers_i/_0638_ ;
 wire \i_ibex/cs_registers_i/_0639_ ;
 wire \i_ibex/cs_registers_i/_0640_ ;
 wire \i_ibex/cs_registers_i/_0641_ ;
 wire \i_ibex/cs_registers_i/_0642_ ;
 wire \i_ibex/cs_registers_i/_0643_ ;
 wire \i_ibex/cs_registers_i/_0644_ ;
 wire \i_ibex/cs_registers_i/_0645_ ;
 wire \i_ibex/cs_registers_i/_0646_ ;
 wire \i_ibex/cs_registers_i/_0647_ ;
 wire \i_ibex/cs_registers_i/_0648_ ;
 wire \i_ibex/cs_registers_i/_0649_ ;
 wire \i_ibex/cs_registers_i/_0650_ ;
 wire \i_ibex/cs_registers_i/_0651_ ;
 wire \i_ibex/cs_registers_i/_0652_ ;
 wire \i_ibex/cs_registers_i/_0653_ ;
 wire \i_ibex/cs_registers_i/_0654_ ;
 wire \i_ibex/cs_registers_i/_0655_ ;
 wire \i_ibex/cs_registers_i/_0656_ ;
 wire \i_ibex/cs_registers_i/_0657_ ;
 wire \i_ibex/cs_registers_i/_0658_ ;
 wire \i_ibex/cs_registers_i/_0659_ ;
 wire \i_ibex/cs_registers_i/_0660_ ;
 wire \i_ibex/cs_registers_i/_0661_ ;
 wire \i_ibex/cs_registers_i/_0662_ ;
 wire \i_ibex/cs_registers_i/_0663_ ;
 wire \i_ibex/cs_registers_i/_0664_ ;
 wire \i_ibex/cs_registers_i/_0665_ ;
 wire net962;
 wire \i_ibex/cs_registers_i/_0667_ ;
 wire \i_ibex/cs_registers_i/_0668_ ;
 wire \i_ibex/cs_registers_i/_0669_ ;
 wire \i_ibex/cs_registers_i/_0670_ ;
 wire \i_ibex/cs_registers_i/_0671_ ;
 wire \i_ibex/cs_registers_i/_0672_ ;
 wire \i_ibex/cs_registers_i/_0673_ ;
 wire \i_ibex/cs_registers_i/_0674_ ;
 wire \i_ibex/cs_registers_i/_0675_ ;
 wire \i_ibex/cs_registers_i/_0676_ ;
 wire \i_ibex/cs_registers_i/_0677_ ;
 wire \i_ibex/cs_registers_i/_0678_ ;
 wire \i_ibex/cs_registers_i/_0679_ ;
 wire \i_ibex/cs_registers_i/_0680_ ;
 wire \i_ibex/cs_registers_i/_0681_ ;
 wire \i_ibex/cs_registers_i/_0682_ ;
 wire \i_ibex/cs_registers_i/_0683_ ;
 wire \i_ibex/cs_registers_i/_0684_ ;
 wire \i_ibex/cs_registers_i/_0685_ ;
 wire \i_ibex/cs_registers_i/_0686_ ;
 wire \i_ibex/cs_registers_i/_0687_ ;
 wire \i_ibex/cs_registers_i/_0688_ ;
 wire \i_ibex/cs_registers_i/_0689_ ;
 wire \i_ibex/cs_registers_i/_0690_ ;
 wire \i_ibex/cs_registers_i/_0691_ ;
 wire \i_ibex/cs_registers_i/_0692_ ;
 wire \i_ibex/cs_registers_i/_0693_ ;
 wire \i_ibex/cs_registers_i/_0694_ ;
 wire \i_ibex/cs_registers_i/_0695_ ;
 wire \i_ibex/cs_registers_i/_0696_ ;
 wire \i_ibex/cs_registers_i/_0697_ ;
 wire \i_ibex/cs_registers_i/_0698_ ;
 wire \i_ibex/cs_registers_i/_0699_ ;
 wire \i_ibex/cs_registers_i/_0700_ ;
 wire \i_ibex/cs_registers_i/_0701_ ;
 wire \i_ibex/cs_registers_i/_0702_ ;
 wire \i_ibex/cs_registers_i/_0703_ ;
 wire \i_ibex/cs_registers_i/_0704_ ;
 wire \i_ibex/cs_registers_i/_0705_ ;
 wire \i_ibex/cs_registers_i/_0706_ ;
 wire \i_ibex/cs_registers_i/_0707_ ;
 wire \i_ibex/cs_registers_i/_0708_ ;
 wire \i_ibex/cs_registers_i/_0709_ ;
 wire \i_ibex/cs_registers_i/_0710_ ;
 wire \i_ibex/cs_registers_i/_0711_ ;
 wire \i_ibex/cs_registers_i/_0712_ ;
 wire \i_ibex/cs_registers_i/_0713_ ;
 wire \i_ibex/cs_registers_i/_0714_ ;
 wire \i_ibex/cs_registers_i/_0715_ ;
 wire \i_ibex/cs_registers_i/_0716_ ;
 wire \i_ibex/cs_registers_i/_0717_ ;
 wire \i_ibex/cs_registers_i/_0718_ ;
 wire \i_ibex/cs_registers_i/_0719_ ;
 wire \i_ibex/cs_registers_i/_0720_ ;
 wire net961;
 wire \i_ibex/cs_registers_i/_0722_ ;
 wire \i_ibex/cs_registers_i/_0723_ ;
 wire \i_ibex/cs_registers_i/_0724_ ;
 wire \i_ibex/cs_registers_i/_0725_ ;
 wire \i_ibex/cs_registers_i/_0726_ ;
 wire \i_ibex/cs_registers_i/_0727_ ;
 wire \i_ibex/cs_registers_i/_0728_ ;
 wire \i_ibex/cs_registers_i/_0729_ ;
 wire \i_ibex/cs_registers_i/_0730_ ;
 wire \i_ibex/cs_registers_i/_0731_ ;
 wire \i_ibex/cs_registers_i/_0732_ ;
 wire \i_ibex/cs_registers_i/_0733_ ;
 wire \i_ibex/cs_registers_i/_0734_ ;
 wire \i_ibex/cs_registers_i/_0735_ ;
 wire \i_ibex/cs_registers_i/_0736_ ;
 wire \i_ibex/cs_registers_i/_0737_ ;
 wire \i_ibex/cs_registers_i/_0738_ ;
 wire \i_ibex/cs_registers_i/_0739_ ;
 wire \i_ibex/cs_registers_i/_0740_ ;
 wire \i_ibex/cs_registers_i/_0741_ ;
 wire \i_ibex/cs_registers_i/_0742_ ;
 wire \i_ibex/cs_registers_i/_0743_ ;
 wire \i_ibex/cs_registers_i/_0744_ ;
 wire \i_ibex/cs_registers_i/_0745_ ;
 wire \i_ibex/cs_registers_i/_0746_ ;
 wire \i_ibex/cs_registers_i/_0747_ ;
 wire \i_ibex/cs_registers_i/_0748_ ;
 wire \i_ibex/cs_registers_i/_0749_ ;
 wire \i_ibex/cs_registers_i/_0750_ ;
 wire \i_ibex/cs_registers_i/_0751_ ;
 wire \i_ibex/cs_registers_i/_0752_ ;
 wire \i_ibex/cs_registers_i/_0753_ ;
 wire \i_ibex/cs_registers_i/_0754_ ;
 wire \i_ibex/cs_registers_i/_0755_ ;
 wire \i_ibex/cs_registers_i/_0756_ ;
 wire \i_ibex/cs_registers_i/_0757_ ;
 wire \i_ibex/cs_registers_i/_0758_ ;
 wire \i_ibex/cs_registers_i/_0759_ ;
 wire \i_ibex/cs_registers_i/_0760_ ;
 wire \i_ibex/cs_registers_i/_0761_ ;
 wire \i_ibex/cs_registers_i/_0762_ ;
 wire \i_ibex/cs_registers_i/_0763_ ;
 wire \i_ibex/cs_registers_i/_0764_ ;
 wire \i_ibex/cs_registers_i/_0765_ ;
 wire \i_ibex/cs_registers_i/_0766_ ;
 wire \i_ibex/cs_registers_i/_0767_ ;
 wire \i_ibex/cs_registers_i/_0768_ ;
 wire \i_ibex/cs_registers_i/_0769_ ;
 wire \i_ibex/cs_registers_i/_0770_ ;
 wire \i_ibex/cs_registers_i/_0771_ ;
 wire \i_ibex/cs_registers_i/_0772_ ;
 wire \i_ibex/cs_registers_i/_0773_ ;
 wire \i_ibex/cs_registers_i/_0774_ ;
 wire \i_ibex/cs_registers_i/_0775_ ;
 wire \i_ibex/cs_registers_i/_0776_ ;
 wire \i_ibex/cs_registers_i/_0777_ ;
 wire \i_ibex/cs_registers_i/_0778_ ;
 wire \i_ibex/cs_registers_i/_0779_ ;
 wire \i_ibex/cs_registers_i/_0780_ ;
 wire \i_ibex/cs_registers_i/_0781_ ;
 wire \i_ibex/cs_registers_i/_0782_ ;
 wire \i_ibex/cs_registers_i/_0783_ ;
 wire \i_ibex/cs_registers_i/_0784_ ;
 wire \i_ibex/cs_registers_i/_0785_ ;
 wire \i_ibex/cs_registers_i/_0786_ ;
 wire \i_ibex/cs_registers_i/_0787_ ;
 wire \i_ibex/cs_registers_i/_0788_ ;
 wire \i_ibex/cs_registers_i/_0789_ ;
 wire \i_ibex/cs_registers_i/_0790_ ;
 wire \i_ibex/cs_registers_i/_0791_ ;
 wire \i_ibex/cs_registers_i/_0792_ ;
 wire \i_ibex/cs_registers_i/_0793_ ;
 wire \i_ibex/cs_registers_i/_0794_ ;
 wire \i_ibex/cs_registers_i/_0795_ ;
 wire \i_ibex/cs_registers_i/_0796_ ;
 wire \i_ibex/cs_registers_i/_0797_ ;
 wire \i_ibex/cs_registers_i/_0798_ ;
 wire \i_ibex/cs_registers_i/_0799_ ;
 wire \i_ibex/cs_registers_i/_0800_ ;
 wire \i_ibex/cs_registers_i/_0801_ ;
 wire \i_ibex/cs_registers_i/_0802_ ;
 wire \i_ibex/cs_registers_i/_0803_ ;
 wire \i_ibex/cs_registers_i/_0804_ ;
 wire \i_ibex/cs_registers_i/_0805_ ;
 wire \i_ibex/cs_registers_i/_0806_ ;
 wire \i_ibex/cs_registers_i/_0807_ ;
 wire \i_ibex/cs_registers_i/_0808_ ;
 wire \i_ibex/cs_registers_i/_0809_ ;
 wire \i_ibex/cs_registers_i/_0810_ ;
 wire \i_ibex/cs_registers_i/_0811_ ;
 wire \i_ibex/cs_registers_i/_0812_ ;
 wire \i_ibex/cs_registers_i/_0813_ ;
 wire \i_ibex/cs_registers_i/_0814_ ;
 wire \i_ibex/cs_registers_i/_0815_ ;
 wire \i_ibex/cs_registers_i/_0816_ ;
 wire \i_ibex/cs_registers_i/_0817_ ;
 wire \i_ibex/cs_registers_i/_0818_ ;
 wire \i_ibex/cs_registers_i/_0819_ ;
 wire \i_ibex/cs_registers_i/_0820_ ;
 wire \i_ibex/cs_registers_i/_0821_ ;
 wire net960;
 wire \i_ibex/cs_registers_i/_0823_ ;
 wire \i_ibex/cs_registers_i/_0824_ ;
 wire \i_ibex/cs_registers_i/_0825_ ;
 wire \i_ibex/cs_registers_i/_0826_ ;
 wire \i_ibex/cs_registers_i/_0827_ ;
 wire \i_ibex/cs_registers_i/_0828_ ;
 wire \i_ibex/cs_registers_i/_0829_ ;
 wire \i_ibex/cs_registers_i/_0830_ ;
 wire \i_ibex/cs_registers_i/_0831_ ;
 wire \i_ibex/cs_registers_i/_0832_ ;
 wire \i_ibex/cs_registers_i/_0833_ ;
 wire \i_ibex/cs_registers_i/_0834_ ;
 wire \i_ibex/cs_registers_i/_0835_ ;
 wire \i_ibex/cs_registers_i/_0836_ ;
 wire \i_ibex/cs_registers_i/_0837_ ;
 wire \i_ibex/cs_registers_i/_0838_ ;
 wire \i_ibex/cs_registers_i/_0839_ ;
 wire \i_ibex/cs_registers_i/_0840_ ;
 wire \i_ibex/cs_registers_i/_0841_ ;
 wire \i_ibex/cs_registers_i/_0842_ ;
 wire \i_ibex/cs_registers_i/_0843_ ;
 wire \i_ibex/cs_registers_i/_0844_ ;
 wire \i_ibex/cs_registers_i/_0845_ ;
 wire \i_ibex/cs_registers_i/_0846_ ;
 wire \i_ibex/cs_registers_i/_0847_ ;
 wire \i_ibex/cs_registers_i/_0848_ ;
 wire \i_ibex/cs_registers_i/_0849_ ;
 wire \i_ibex/cs_registers_i/_0850_ ;
 wire \i_ibex/cs_registers_i/_0851_ ;
 wire \i_ibex/cs_registers_i/_0852_ ;
 wire \i_ibex/cs_registers_i/_0853_ ;
 wire \i_ibex/cs_registers_i/_0854_ ;
 wire \i_ibex/cs_registers_i/_0855_ ;
 wire \i_ibex/cs_registers_i/_0856_ ;
 wire \i_ibex/cs_registers_i/_0857_ ;
 wire \i_ibex/cs_registers_i/_0858_ ;
 wire \i_ibex/cs_registers_i/_0859_ ;
 wire \i_ibex/cs_registers_i/_0860_ ;
 wire \i_ibex/cs_registers_i/_0861_ ;
 wire \i_ibex/cs_registers_i/_0862_ ;
 wire \i_ibex/cs_registers_i/_0863_ ;
 wire \i_ibex/cs_registers_i/_0864_ ;
 wire net959;
 wire \i_ibex/cs_registers_i/_0866_ ;
 wire net958;
 wire \i_ibex/cs_registers_i/_0868_ ;
 wire net957;
 wire \i_ibex/cs_registers_i/_0870_ ;
 wire net956;
 wire net955;
 wire \i_ibex/cs_registers_i/_0873_ ;
 wire net954;
 wire net953;
 wire \i_ibex/cs_registers_i/_0876_ ;
 wire \i_ibex/cs_registers_i/_0877_ ;
 wire \i_ibex/cs_registers_i/_0878_ ;
 wire \i_ibex/cs_registers_i/_0879_ ;
 wire \i_ibex/cs_registers_i/_0880_ ;
 wire \i_ibex/cs_registers_i/_0881_ ;
 wire net952;
 wire net951;
 wire \i_ibex/cs_registers_i/_0884_ ;
 wire net950;
 wire \i_ibex/cs_registers_i/_0886_ ;
 wire \i_ibex/cs_registers_i/_0887_ ;
 wire \i_ibex/cs_registers_i/_0888_ ;
 wire \i_ibex/cs_registers_i/_0889_ ;
 wire net949;
 wire \i_ibex/cs_registers_i/_0891_ ;
 wire \i_ibex/cs_registers_i/_0892_ ;
 wire net948;
 wire \i_ibex/cs_registers_i/_0894_ ;
 wire \i_ibex/cs_registers_i/_0895_ ;
 wire \i_ibex/cs_registers_i/_0896_ ;
 wire \i_ibex/cs_registers_i/_0897_ ;
 wire \i_ibex/cs_registers_i/_0898_ ;
 wire \i_ibex/cs_registers_i/_0899_ ;
 wire \i_ibex/cs_registers_i/_0900_ ;
 wire \i_ibex/cs_registers_i/_0901_ ;
 wire \i_ibex/cs_registers_i/_0902_ ;
 wire \i_ibex/cs_registers_i/_0903_ ;
 wire \i_ibex/cs_registers_i/_0904_ ;
 wire \i_ibex/cs_registers_i/_0905_ ;
 wire net947;
 wire \i_ibex/cs_registers_i/_0907_ ;
 wire \i_ibex/cs_registers_i/_0908_ ;
 wire \i_ibex/cs_registers_i/_0909_ ;
 wire \i_ibex/cs_registers_i/_0910_ ;
 wire \i_ibex/cs_registers_i/_0911_ ;
 wire \i_ibex/cs_registers_i/_0912_ ;
 wire \i_ibex/cs_registers_i/_0913_ ;
 wire \i_ibex/cs_registers_i/_0914_ ;
 wire \i_ibex/cs_registers_i/_0915_ ;
 wire \i_ibex/cs_registers_i/_0916_ ;
 wire \i_ibex/cs_registers_i/_0917_ ;
 wire \i_ibex/cs_registers_i/_0918_ ;
 wire \i_ibex/cs_registers_i/_0919_ ;
 wire \i_ibex/cs_registers_i/_0920_ ;
 wire \i_ibex/cs_registers_i/_0921_ ;
 wire \i_ibex/cs_registers_i/_0922_ ;
 wire \i_ibex/cs_registers_i/_0923_ ;
 wire \i_ibex/cs_registers_i/_0924_ ;
 wire \i_ibex/cs_registers_i/_0925_ ;
 wire \i_ibex/cs_registers_i/_0926_ ;
 wire \i_ibex/cs_registers_i/_0927_ ;
 wire \i_ibex/cs_registers_i/_0928_ ;
 wire \i_ibex/cs_registers_i/_0929_ ;
 wire \i_ibex/cs_registers_i/_0930_ ;
 wire \i_ibex/cs_registers_i/_0931_ ;
 wire \i_ibex/cs_registers_i/_0932_ ;
 wire \i_ibex/cs_registers_i/_0933_ ;
 wire \i_ibex/cs_registers_i/_0934_ ;
 wire \i_ibex/cs_registers_i/_0935_ ;
 wire \i_ibex/cs_registers_i/_0936_ ;
 wire \i_ibex/cs_registers_i/_0937_ ;
 wire \i_ibex/cs_registers_i/_0938_ ;
 wire \i_ibex/cs_registers_i/_0939_ ;
 wire \i_ibex/cs_registers_i/_0940_ ;
 wire \i_ibex/cs_registers_i/_0941_ ;
 wire \i_ibex/cs_registers_i/_0942_ ;
 wire \i_ibex/cs_registers_i/_0943_ ;
 wire \i_ibex/cs_registers_i/_0944_ ;
 wire \i_ibex/cs_registers_i/_0945_ ;
 wire net946;
 wire \i_ibex/cs_registers_i/_0947_ ;
 wire \i_ibex/cs_registers_i/_0948_ ;
 wire net945;
 wire \i_ibex/cs_registers_i/_0950_ ;
 wire net944;
 wire \i_ibex/cs_registers_i/_0952_ ;
 wire net943;
 wire \i_ibex/cs_registers_i/_0954_ ;
 wire \i_ibex/cs_registers_i/_0955_ ;
 wire \i_ibex/cs_registers_i/_0956_ ;
 wire net942;
 wire net941;
 wire \i_ibex/cs_registers_i/_0959_ ;
 wire \i_ibex/cs_registers_i/_0960_ ;
 wire \i_ibex/cs_registers_i/_0961_ ;
 wire \i_ibex/cs_registers_i/_0962_ ;
 wire \i_ibex/cs_registers_i/_0963_ ;
 wire \i_ibex/cs_registers_i/_0964_ ;
 wire \i_ibex/cs_registers_i/_0965_ ;
 wire net940;
 wire \i_ibex/cs_registers_i/_0967_ ;
 wire \i_ibex/cs_registers_i/_0968_ ;
 wire \i_ibex/cs_registers_i/_0969_ ;
 wire \i_ibex/cs_registers_i/_0970_ ;
 wire \i_ibex/cs_registers_i/_0971_ ;
 wire \i_ibex/cs_registers_i/_0972_ ;
 wire \i_ibex/cs_registers_i/_0973_ ;
 wire \i_ibex/cs_registers_i/_0974_ ;
 wire \i_ibex/cs_registers_i/_0975_ ;
 wire \i_ibex/cs_registers_i/_0976_ ;
 wire \i_ibex/cs_registers_i/_0977_ ;
 wire net938;
 wire \i_ibex/cs_registers_i/_0979_ ;
 wire \i_ibex/cs_registers_i/_0980_ ;
 wire \i_ibex/cs_registers_i/_0981_ ;
 wire \i_ibex/cs_registers_i/_0982_ ;
 wire \i_ibex/cs_registers_i/_0983_ ;
 wire \i_ibex/cs_registers_i/_0984_ ;
 wire net937;
 wire \i_ibex/cs_registers_i/_0986_ ;
 wire \i_ibex/cs_registers_i/_0987_ ;
 wire \i_ibex/cs_registers_i/_0988_ ;
 wire \i_ibex/cs_registers_i/_0989_ ;
 wire \i_ibex/cs_registers_i/_0990_ ;
 wire \i_ibex/cs_registers_i/_0991_ ;
 wire net936;
 wire \i_ibex/cs_registers_i/_0993_ ;
 wire \i_ibex/cs_registers_i/_0994_ ;
 wire \i_ibex/cs_registers_i/_0995_ ;
 wire \i_ibex/cs_registers_i/_0996_ ;
 wire \i_ibex/cs_registers_i/_0997_ ;
 wire \i_ibex/cs_registers_i/_0998_ ;
 wire \i_ibex/cs_registers_i/_0999_ ;
 wire \i_ibex/cs_registers_i/_1000_ ;
 wire \i_ibex/cs_registers_i/_1001_ ;
 wire \i_ibex/cs_registers_i/_1002_ ;
 wire \i_ibex/cs_registers_i/_1003_ ;
 wire \i_ibex/cs_registers_i/_1004_ ;
 wire \i_ibex/cs_registers_i/_1005_ ;
 wire \i_ibex/cs_registers_i/_1006_ ;
 wire \i_ibex/cs_registers_i/_1007_ ;
 wire \i_ibex/cs_registers_i/_1008_ ;
 wire \i_ibex/cs_registers_i/_1009_ ;
 wire \i_ibex/cs_registers_i/_1010_ ;
 wire \i_ibex/cs_registers_i/_1011_ ;
 wire \i_ibex/cs_registers_i/_1012_ ;
 wire \i_ibex/cs_registers_i/_1013_ ;
 wire \i_ibex/cs_registers_i/_1014_ ;
 wire \i_ibex/cs_registers_i/_1015_ ;
 wire \i_ibex/cs_registers_i/_1016_ ;
 wire \i_ibex/cs_registers_i/_1017_ ;
 wire \i_ibex/cs_registers_i/_1018_ ;
 wire \i_ibex/cs_registers_i/_1019_ ;
 wire \i_ibex/cs_registers_i/_1020_ ;
 wire \i_ibex/cs_registers_i/_1021_ ;
 wire \i_ibex/cs_registers_i/_1022_ ;
 wire \i_ibex/cs_registers_i/_1023_ ;
 wire \i_ibex/cs_registers_i/_1024_ ;
 wire \i_ibex/cs_registers_i/_1025_ ;
 wire \i_ibex/cs_registers_i/_1026_ ;
 wire \i_ibex/cs_registers_i/_1027_ ;
 wire \i_ibex/cs_registers_i/_1028_ ;
 wire \i_ibex/cs_registers_i/_1029_ ;
 wire \i_ibex/cs_registers_i/_1030_ ;
 wire \i_ibex/cs_registers_i/_1031_ ;
 wire \i_ibex/cs_registers_i/_1032_ ;
 wire \i_ibex/cs_registers_i/_1033_ ;
 wire \i_ibex/cs_registers_i/_1034_ ;
 wire \i_ibex/cs_registers_i/_1035_ ;
 wire \i_ibex/cs_registers_i/_1036_ ;
 wire \i_ibex/cs_registers_i/_1037_ ;
 wire \i_ibex/cs_registers_i/_1038_ ;
 wire \i_ibex/cs_registers_i/_1039_ ;
 wire \i_ibex/cs_registers_i/_1040_ ;
 wire \i_ibex/cs_registers_i/_1041_ ;
 wire \i_ibex/cs_registers_i/_1042_ ;
 wire \i_ibex/cs_registers_i/_1043_ ;
 wire \i_ibex/cs_registers_i/_1044_ ;
 wire \i_ibex/cs_registers_i/_1045_ ;
 wire \i_ibex/cs_registers_i/_1046_ ;
 wire \i_ibex/cs_registers_i/_1047_ ;
 wire \i_ibex/cs_registers_i/_1048_ ;
 wire \i_ibex/cs_registers_i/_1049_ ;
 wire \i_ibex/cs_registers_i/_1050_ ;
 wire \i_ibex/cs_registers_i/_1051_ ;
 wire \i_ibex/cs_registers_i/_1052_ ;
 wire \i_ibex/cs_registers_i/_1053_ ;
 wire \i_ibex/cs_registers_i/_1054_ ;
 wire \i_ibex/cs_registers_i/_1055_ ;
 wire \i_ibex/cs_registers_i/_1056_ ;
 wire \i_ibex/cs_registers_i/_1057_ ;
 wire \i_ibex/cs_registers_i/_1058_ ;
 wire \i_ibex/cs_registers_i/_1059_ ;
 wire \i_ibex/cs_registers_i/_1060_ ;
 wire \i_ibex/cs_registers_i/_1061_ ;
 wire \i_ibex/cs_registers_i/_1062_ ;
 wire \i_ibex/cs_registers_i/_1063_ ;
 wire \i_ibex/cs_registers_i/_1064_ ;
 wire \i_ibex/cs_registers_i/_1065_ ;
 wire \i_ibex/cs_registers_i/_1066_ ;
 wire \i_ibex/cs_registers_i/_1067_ ;
 wire \i_ibex/cs_registers_i/_1068_ ;
 wire \i_ibex/cs_registers_i/_1069_ ;
 wire \i_ibex/cs_registers_i/_1070_ ;
 wire \i_ibex/cs_registers_i/_1071_ ;
 wire net935;
 wire net934;
 wire net933;
 wire \i_ibex/cs_registers_i/_1075_ ;
 wire net932;
 wire \i_ibex/cs_registers_i/_1077_ ;
 wire \i_ibex/cs_registers_i/_1078_ ;
 wire net931;
 wire net930;
 wire net929;
 wire \i_ibex/cs_registers_i/_1082_ ;
 wire \i_ibex/cs_registers_i/_1083_ ;
 wire \i_ibex/cs_registers_i/_1084_ ;
 wire \i_ibex/cs_registers_i/_1085_ ;
 wire \i_ibex/cs_registers_i/_1086_ ;
 wire \i_ibex/cs_registers_i/_1087_ ;
 wire \i_ibex/cs_registers_i/_1088_ ;
 wire \i_ibex/cs_registers_i/_1089_ ;
 wire \i_ibex/cs_registers_i/_1090_ ;
 wire \i_ibex/cs_registers_i/_1091_ ;
 wire \i_ibex/cs_registers_i/_1092_ ;
 wire \i_ibex/cs_registers_i/_1093_ ;
 wire \i_ibex/cs_registers_i/_1094_ ;
 wire \i_ibex/cs_registers_i/_1095_ ;
 wire \i_ibex/cs_registers_i/_1096_ ;
 wire \i_ibex/cs_registers_i/_1097_ ;
 wire \i_ibex/cs_registers_i/_1098_ ;
 wire \i_ibex/cs_registers_i/_1099_ ;
 wire \i_ibex/cs_registers_i/_1100_ ;
 wire \i_ibex/cs_registers_i/_1101_ ;
 wire \i_ibex/cs_registers_i/_1102_ ;
 wire \i_ibex/cs_registers_i/_1103_ ;
 wire \i_ibex/cs_registers_i/_1104_ ;
 wire \i_ibex/cs_registers_i/_1105_ ;
 wire \i_ibex/cs_registers_i/_1106_ ;
 wire \i_ibex/cs_registers_i/_1107_ ;
 wire \i_ibex/cs_registers_i/_1108_ ;
 wire \i_ibex/cs_registers_i/_1109_ ;
 wire \i_ibex/cs_registers_i/_1110_ ;
 wire \i_ibex/cs_registers_i/_1111_ ;
 wire \i_ibex/cs_registers_i/_1112_ ;
 wire \i_ibex/cs_registers_i/_1113_ ;
 wire \i_ibex/cs_registers_i/_1114_ ;
 wire \i_ibex/cs_registers_i/_1115_ ;
 wire \i_ibex/cs_registers_i/_1116_ ;
 wire \i_ibex/cs_registers_i/_1117_ ;
 wire \i_ibex/cs_registers_i/_1118_ ;
 wire \i_ibex/cs_registers_i/_1119_ ;
 wire \i_ibex/cs_registers_i/_1120_ ;
 wire \i_ibex/cs_registers_i/_1121_ ;
 wire \i_ibex/cs_registers_i/_1122_ ;
 wire \i_ibex/cs_registers_i/_1123_ ;
 wire \i_ibex/cs_registers_i/_1124_ ;
 wire \i_ibex/cs_registers_i/_1125_ ;
 wire \i_ibex/cs_registers_i/_1126_ ;
 wire \i_ibex/cs_registers_i/_1127_ ;
 wire net1049;
 wire \i_ibex/cs_registers_i/dcsr_en ;
 wire \i_ibex/cs_registers_i/depc_en ;
 wire \i_ibex/cs_registers_i/dscratch0_en ;
 wire \i_ibex/cs_registers_i/dscratch1_en ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_control ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.tmatch_control_we ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.tmatch_value_we ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.tselect_q ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.tselect_we ;
 wire \i_ibex/cs_registers_i/instr_ret_i_$_AND__A_B ;
 wire \i_ibex/cs_registers_i/mcause_en ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ;
 wire \i_ibex/cs_registers_i/mepc_en ;
 wire \i_ibex/cs_registers_i/mie_en ;
 wire \i_ibex/cs_registers_i/minstret_counter_i_counter_inc_i ;
 wire \i_ibex/cs_registers_i/mscratch_en ;
 wire net939;
 wire \i_ibex/cs_registers_i/mstatus_en ;
 wire \i_ibex/cs_registers_i/mtval_en ;
 wire \i_ibex/cs_registers_i/mtvec_en ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/_0_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/_1_ ;
 wire net71;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_000_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_001_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_002_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_003_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_004_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_005_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_006_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_007_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_008_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_009_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_010_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_011_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_012_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_013_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_014_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_015_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_016_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_017_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_018_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_019_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_020_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_021_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_022_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_023_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_024_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_025_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_026_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_027_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_028_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_029_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_030_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_031_ ;
 wire net926;
 wire net925;
 wire net928;
 wire net927;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_036_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_037_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_038_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_039_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_040_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_041_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_042_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_043_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_044_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_045_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_046_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_047_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_048_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_049_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_050_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_051_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_052_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_053_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_054_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_055_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_056_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_057_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_058_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_059_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_060_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_061_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_062_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_063_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_064_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_065_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_066_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_067_ ;
 wire net70;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_0_ ;
 wire \i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_1_ ;
 wire net69;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_000_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_001_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_002_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_003_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_004_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_005_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_006_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_007_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_008_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_009_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_010_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_011_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_012_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_013_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_014_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_015_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_016_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_017_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_018_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_019_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_020_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_021_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_022_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_023_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_024_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_025_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_026_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_027_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_028_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_029_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_030_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_031_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_032_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_033_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_034_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_035_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_036_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_037_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_038_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_039_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_040_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_041_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_042_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_043_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_044_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_045_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_046_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_047_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_048_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_049_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_050_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_051_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_052_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_053_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_054_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_055_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_056_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_057_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_058_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_059_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_060_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_061_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_062_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_063_ ;
 wire net924;
 wire net923;
 wire net922;
 wire net921;
 wire net920;
 wire net919;
 wire net918;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_071_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_072_ ;
 wire net917;
 wire net916;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_075_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_076_ ;
 wire net915;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_078_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_079_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_080_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_081_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_082_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_083_ ;
 wire net914;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_085_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_086_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_087_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_088_ ;
 wire net913;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_090_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_091_ ;
 wire net912;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_093_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_094_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_095_ ;
 wire net911;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_097_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_098_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_099_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_100_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_101_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_102_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_103_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_104_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_105_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_106_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_107_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_108_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_109_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_110_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_111_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_112_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_113_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_114_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_115_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_116_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_117_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_118_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_119_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_120_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_121_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_122_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_123_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_124_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_125_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_126_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_127_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_128_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_129_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_130_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_131_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_132_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_133_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_134_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_135_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_136_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_137_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_138_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_139_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_140_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_141_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_142_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_143_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_144_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_145_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_146_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_147_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_148_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_149_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_150_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_151_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_152_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_153_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_154_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_155_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_156_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_157_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_158_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_159_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_160_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_161_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_162_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_163_ ;
 wire net910;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_165_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_166_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_167_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_168_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_169_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_170_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_171_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_172_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_173_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_174_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_175_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_176_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_177_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_178_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_179_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_180_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_181_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_182_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_183_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_184_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_185_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_186_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_187_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_188_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_189_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_190_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_191_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_192_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_193_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_194_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_195_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_196_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_197_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_198_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_199_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_200_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_201_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_202_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_203_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_204_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_205_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_206_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_207_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_208_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_209_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_210_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_211_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_212_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_213_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_214_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_215_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_216_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_217_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_218_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_219_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_220_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_221_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_222_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_223_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_224_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_225_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_226_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_227_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_228_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_229_ ;
 wire net909;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_231_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_232_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_233_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_234_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_235_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_236_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_237_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_238_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_239_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_240_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_241_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_242_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_243_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_244_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_245_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_246_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_247_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_248_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_249_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_250_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_251_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_252_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_253_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_254_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_255_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_256_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_257_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_258_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_259_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_260_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_261_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_262_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_263_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_264_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_265_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_266_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_267_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_268_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_269_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_270_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_271_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_272_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_273_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_274_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_275_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_276_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_277_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_278_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_279_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_280_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_281_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_282_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_283_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_284_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_285_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_286_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_287_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_288_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_289_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_290_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_291_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_292_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_293_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_294_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_295_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_296_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_297_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_298_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_299_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_300_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_301_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_302_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_303_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_304_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_305_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_306_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_307_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_308_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_309_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_310_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_311_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_312_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_313_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_314_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_315_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_316_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_317_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_318_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_319_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_320_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_321_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_322_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_323_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_324_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_325_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_326_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_327_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_328_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_329_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_330_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_331_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_332_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_333_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_334_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_335_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_336_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_337_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_338_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_339_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_340_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_341_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_342_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_343_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_344_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_345_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_346_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_347_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_348_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_349_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_350_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_351_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_352_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_353_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_354_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_355_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_356_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_357_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_358_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_359_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_360_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_361_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_362_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_363_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_364_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_365_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_366_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_367_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_368_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_369_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_370_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_371_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_372_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_373_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_374_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_375_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_376_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_377_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_378_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_379_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_380_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_381_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_382_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_383_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_384_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_385_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_386_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_387_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_388_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_389_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_390_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_391_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_392_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_393_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_394_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_395_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_396_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_397_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_398_ ;
 wire \i_ibex/cs_registers_i/mcycle_counter_i/_399_ ;
 wire net68;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0000_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0001_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0002_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0003_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0004_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0005_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0006_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0007_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0008_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0009_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0010_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0011_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0012_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0013_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0014_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0015_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0016_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0017_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0018_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0019_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0020_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0021_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0022_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0023_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0024_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0025_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0026_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0027_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0028_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0029_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0030_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0031_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0032_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0033_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0034_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0035_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0036_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0037_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0038_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0039_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0040_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0041_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0042_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0043_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0044_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0045_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0046_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0047_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0048_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0049_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0050_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0051_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0052_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0053_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0054_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0055_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0056_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0057_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0058_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0059_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0060_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0061_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0062_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0063_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0064_ ;
 wire net908;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0066_ ;
 wire net907;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0068_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0069_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0070_ ;
 wire net906;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0072_ ;
 wire net905;
 wire net904;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0075_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0076_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0077_ ;
 wire net903;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0079_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0080_ ;
 wire net902;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0082_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0083_ ;
 wire net901;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0085_ ;
 wire net900;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0087_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0088_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0089_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0090_ ;
 wire net899;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0092_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0093_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0094_ ;
 wire net898;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0096_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0097_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0098_ ;
 wire net897;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0100_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0101_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0102_ ;
 wire net896;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0104_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0105_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0106_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0107_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0108_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0109_ ;
 wire net895;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0111_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0112_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0113_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0114_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0115_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0116_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0117_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0118_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0119_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0120_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0121_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0122_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0123_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0124_ ;
 wire net894;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0126_ ;
 wire net893;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0128_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0129_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0130_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0131_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0132_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0133_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0134_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0135_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0136_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0137_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0138_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0139_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0140_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0141_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0142_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0143_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0144_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0145_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0146_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0147_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0148_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0149_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0150_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0151_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0152_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0153_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0154_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0155_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0156_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0157_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0158_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0159_ ;
 wire net892;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0161_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0162_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0163_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0164_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0165_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0166_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0167_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0168_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0169_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0170_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0171_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0172_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0173_ ;
 wire net891;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0175_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0176_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0177_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0178_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0179_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0180_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0181_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0182_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0183_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0184_ ;
 wire net890;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0186_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0187_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0188_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0189_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0190_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0191_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0192_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0193_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0194_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0195_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0196_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0197_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0198_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0199_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0200_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0201_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0202_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0203_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0204_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0205_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0206_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0207_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0208_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0209_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0210_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0211_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0212_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0213_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0214_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0215_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0216_ ;
 wire net889;
 wire net888;
 wire net887;
 wire net886;
 wire net885;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0222_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0223_ ;
 wire net884;
 wire net883;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0226_ ;
 wire net882;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0228_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0229_ ;
 wire net881;
 wire net880;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0232_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0233_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0234_ ;
 wire net879;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0236_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0237_ ;
 wire net878;
 wire net877;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0240_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0241_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0242_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0243_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0244_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0245_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0246_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0247_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0248_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0249_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0250_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0251_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0252_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0253_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0254_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0255_ ;
 wire net876;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0257_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0258_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0259_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0260_ ;
 wire net875;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0262_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0263_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0264_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0265_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0266_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0267_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0268_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0269_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0270_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0271_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0272_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0273_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0274_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0275_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0276_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0277_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0278_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0279_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0280_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0281_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0282_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0283_ ;
 wire net874;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0285_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0286_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0287_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0288_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0289_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0290_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0291_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0292_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0293_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0294_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0295_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0296_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0297_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0298_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0299_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0300_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0301_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0302_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0303_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0304_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0305_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0306_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0307_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0308_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0309_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0310_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0311_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0312_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0313_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0314_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0315_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0316_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0317_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0318_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0319_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0320_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0321_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0322_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0323_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0324_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0325_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0326_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0327_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0328_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0329_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0330_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0331_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0332_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0333_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0334_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0335_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0336_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0337_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0338_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0339_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0340_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0341_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0342_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0343_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0344_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0345_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0346_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0347_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0348_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0349_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0350_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0351_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0352_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0353_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0354_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0355_ ;
 wire net873;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0357_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0358_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0359_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0360_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0361_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0362_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0363_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0364_ ;
 wire net872;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0366_ ;
 wire net871;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0368_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0369_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0370_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0371_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0372_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0373_ ;
 wire net870;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0375_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0376_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0377_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0378_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0379_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0380_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0381_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0382_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0383_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0384_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0385_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0386_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0387_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0388_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0389_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0390_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0391_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0392_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0393_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0394_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0395_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0396_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0397_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0398_ ;
 wire net869;
 wire net868;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0401_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0402_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0403_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0404_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0405_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0406_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0407_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0408_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0409_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0410_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0411_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0412_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0413_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0414_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0415_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0416_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0417_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0418_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0419_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0420_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0421_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0422_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0423_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0424_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0425_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0426_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0427_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0428_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0429_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0430_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0431_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0432_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0433_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0434_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0435_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0436_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0437_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0438_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0439_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0440_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0441_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0442_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0443_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0444_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0445_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0446_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0447_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0448_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0449_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0450_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0451_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0452_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0453_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0454_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0455_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0456_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0457_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0458_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0459_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0460_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0461_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0462_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0463_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0464_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0465_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0466_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0467_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0468_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0469_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0470_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0471_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0472_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0473_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0474_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0475_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0476_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0477_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0478_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0479_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0480_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0481_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0482_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0483_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0484_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0485_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0486_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0487_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0488_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0489_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0490_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0491_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0492_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0493_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0494_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0495_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0496_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0497_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0498_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0499_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0500_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0501_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0502_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0503_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0504_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0505_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0506_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0507_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0508_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0509_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0510_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0511_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0512_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0513_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0514_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0515_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0516_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0517_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0518_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0519_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0520_ ;
 wire \i_ibex/cs_registers_i/minstret_counter_i/_0521_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_031_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_032_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_033_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_034_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_035_ ;
 wire net865;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_037_ ;
 wire net864;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_039_ ;
 wire net867;
 wire net866;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_067_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_068_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_069_ ;
 wire \i_ibex/cs_registers_i/u_dcsr_csr/_070_ ;
 wire net67;
 wire \i_ibex/cs_registers_i/u_depc_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_031_ ;
 wire net861;
 wire net860;
 wire net863;
 wire net862;
 wire \i_ibex/cs_registers_i/u_depc_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_depc_csr/_067_ ;
 wire net66;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_031_ ;
 wire net857;
 wire net856;
 wire net859;
 wire net858;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_dscratch0_csr/_067_ ;
 wire net65;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_031_ ;
 wire net853;
 wire net852;
 wire net855;
 wire net854;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_dscratch1_csr/_067_ ;
 wire net64;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_00_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_01_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_02_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_03_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_04_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_05_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_06_ ;
 wire net851;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_08_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_09_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_10_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_11_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_12_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_13_ ;
 wire \i_ibex/cs_registers_i/u_mcause_csr/_14_ ;
 wire net63;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_031_ ;
 wire net848;
 wire net847;
 wire net850;
 wire net849;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_mepc_csr/_067_ ;
 wire net62;
 wire \i_ibex/cs_registers_i/u_mie_csr/_00_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_01_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_02_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_03_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_04_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_05_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_06_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_07_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_08_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_09_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_10_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_11_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_12_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_13_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_14_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_15_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_16_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_17_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_18_ ;
 wire net846;
 wire net845;
 wire \i_ibex/cs_registers_i/u_mie_csr/_21_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_22_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_23_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_24_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_25_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_26_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_27_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_28_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_29_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_30_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_31_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_32_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_33_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_34_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_35_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_36_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_37_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_38_ ;
 wire \i_ibex/cs_registers_i/u_mie_csr/_39_ ;
 wire net61;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_031_ ;
 wire net842;
 wire net841;
 wire net844;
 wire net843;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_mscratch_csr/_067_ ;
 wire net60;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_00_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_01_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_02_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_03_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_04_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_05_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_06_ ;
 wire net840;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_08_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_09_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_10_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_11_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_12_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_13_ ;
 wire \i_ibex/cs_registers_i/u_mstack_cause_csr/_14_ ;
 wire net59;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_00_ ;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_01_ ;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_02_ ;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_03_ ;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_04_ ;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_05_ ;
 wire \i_ibex/cs_registers_i/u_mstack_csr/_06_ ;
 wire net58;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_031_ ;
 wire net837;
 wire net836;
 wire net839;
 wire net838;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_mstack_epc_csr/_067_ ;
 wire net57;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_00_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_01_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_02_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_03_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_04_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_05_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_06_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_07_ ;
 wire net835;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_09_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_10_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_11_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_12_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_13_ ;
 wire \i_ibex/cs_registers_i/u_mstatus_csr/_14_ ;
 wire net56;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_031_ ;
 wire net832;
 wire net831;
 wire net834;
 wire net833;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_036_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_037_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_mtval_csr/_067_ ;
 wire net55;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_000_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_001_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_002_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_003_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_004_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_005_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_006_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_007_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_008_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_009_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_010_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_011_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_012_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_013_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_014_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_015_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_016_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_017_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_018_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_019_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_020_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_021_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_022_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_023_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_024_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_025_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_026_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_027_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_028_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_029_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_030_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_031_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_032_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_033_ ;
 wire net828;
 wire net827;
 wire net830;
 wire net829;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_038_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_039_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_040_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_041_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_042_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_043_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_044_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_045_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_046_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_047_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_048_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_049_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_050_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_051_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_052_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_053_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_054_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_055_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_056_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_057_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_058_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_059_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_060_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_061_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_062_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_063_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_064_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_065_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_066_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_067_ ;
 wire \i_ibex/cs_registers_i/u_mtvec_csr/_068_ ;
 wire net54;
 wire \i_ibex/ex_block_i/alu_is_equal_result ;
 wire \i_ibex/ex_block_i/alu_i/_0000_ ;
 wire \i_ibex/ex_block_i/alu_i/_0001_ ;
 wire \i_ibex/ex_block_i/alu_i/_0002_ ;
 wire \i_ibex/ex_block_i/alu_i/_0003_ ;
 wire \i_ibex/ex_block_i/alu_i/_0004_ ;
 wire \i_ibex/ex_block_i/alu_i/_0005_ ;
 wire \i_ibex/ex_block_i/alu_i/_0006_ ;
 wire \i_ibex/ex_block_i/alu_i/_0007_ ;
 wire \i_ibex/ex_block_i/alu_i/_0008_ ;
 wire \i_ibex/ex_block_i/alu_i/_0009_ ;
 wire \i_ibex/ex_block_i/alu_i/_0010_ ;
 wire \i_ibex/ex_block_i/alu_i/_0011_ ;
 wire \i_ibex/ex_block_i/alu_i/_0012_ ;
 wire \i_ibex/ex_block_i/alu_i/_0013_ ;
 wire \i_ibex/ex_block_i/alu_i/_0014_ ;
 wire \i_ibex/ex_block_i/alu_i/_0015_ ;
 wire \i_ibex/ex_block_i/alu_i/_0016_ ;
 wire \i_ibex/ex_block_i/alu_i/_0017_ ;
 wire \i_ibex/ex_block_i/alu_i/_0018_ ;
 wire \i_ibex/ex_block_i/alu_i/_0019_ ;
 wire \i_ibex/ex_block_i/alu_i/_0020_ ;
 wire \i_ibex/ex_block_i/alu_i/_0021_ ;
 wire \i_ibex/ex_block_i/alu_i/_0022_ ;
 wire \i_ibex/ex_block_i/alu_i/_0023_ ;
 wire \i_ibex/ex_block_i/alu_i/_0024_ ;
 wire \i_ibex/ex_block_i/alu_i/_0025_ ;
 wire \i_ibex/ex_block_i/alu_i/_0026_ ;
 wire \i_ibex/ex_block_i/alu_i/_0027_ ;
 wire \i_ibex/ex_block_i/alu_i/_0028_ ;
 wire \i_ibex/ex_block_i/alu_i/_0029_ ;
 wire \i_ibex/ex_block_i/alu_i/_0030_ ;
 wire \i_ibex/ex_block_i/alu_i/_0031_ ;
 wire \i_ibex/ex_block_i/alu_i/_0032_ ;
 wire \i_ibex/ex_block_i/alu_i/_0033_ ;
 wire \i_ibex/ex_block_i/alu_i/_0034_ ;
 wire \i_ibex/ex_block_i/alu_i/_0035_ ;
 wire \i_ibex/ex_block_i/alu_i/_0036_ ;
 wire \i_ibex/ex_block_i/alu_i/_0037_ ;
 wire \i_ibex/ex_block_i/alu_i/_0038_ ;
 wire \i_ibex/ex_block_i/alu_i/_0039_ ;
 wire \i_ibex/ex_block_i/alu_i/_0040_ ;
 wire \i_ibex/ex_block_i/alu_i/_0041_ ;
 wire \i_ibex/ex_block_i/alu_i/_0042_ ;
 wire \i_ibex/ex_block_i/alu_i/_0043_ ;
 wire \i_ibex/ex_block_i/alu_i/_0044_ ;
 wire \i_ibex/ex_block_i/alu_i/_0045_ ;
 wire \i_ibex/ex_block_i/alu_i/_0046_ ;
 wire \i_ibex/ex_block_i/alu_i/_0047_ ;
 wire \i_ibex/ex_block_i/alu_i/_0048_ ;
 wire \i_ibex/ex_block_i/alu_i/_0049_ ;
 wire \i_ibex/ex_block_i/alu_i/_0050_ ;
 wire \i_ibex/ex_block_i/alu_i/_0051_ ;
 wire \i_ibex/ex_block_i/alu_i/_0052_ ;
 wire \i_ibex/ex_block_i/alu_i/_0053_ ;
 wire \i_ibex/ex_block_i/alu_i/_0054_ ;
 wire \i_ibex/ex_block_i/alu_i/_0055_ ;
 wire \i_ibex/ex_block_i/alu_i/_0056_ ;
 wire \i_ibex/ex_block_i/alu_i/_0057_ ;
 wire \i_ibex/ex_block_i/alu_i/_0058_ ;
 wire \i_ibex/ex_block_i/alu_i/_0059_ ;
 wire \i_ibex/ex_block_i/alu_i/_0060_ ;
 wire \i_ibex/ex_block_i/alu_i/_0061_ ;
 wire \i_ibex/ex_block_i/alu_i/_0062_ ;
 wire \i_ibex/ex_block_i/alu_i/_0063_ ;
 wire \i_ibex/ex_block_i/alu_i/_0064_ ;
 wire \i_ibex/ex_block_i/alu_i/_0065_ ;
 wire \i_ibex/ex_block_i/alu_i/_0066_ ;
 wire \i_ibex/ex_block_i/alu_i/_0067_ ;
 wire \i_ibex/ex_block_i/alu_i/_0068_ ;
 wire \i_ibex/ex_block_i/alu_i/_0069_ ;
 wire \i_ibex/ex_block_i/alu_i/_0070_ ;
 wire \i_ibex/ex_block_i/alu_i/_0071_ ;
 wire \i_ibex/ex_block_i/alu_i/_0072_ ;
 wire net744;
 wire net743;
 wire net742;
 wire \i_ibex/ex_block_i/alu_i/_0076_ ;
 wire net741;
 wire net740;
 wire net739;
 wire net738;
 wire \i_ibex/ex_block_i/alu_i/_0081_ ;
 wire \i_ibex/ex_block_i/alu_i/_0082_ ;
 wire \i_ibex/ex_block_i/alu_i/_0083_ ;
 wire net737;
 wire \i_ibex/ex_block_i/alu_i/_0085_ ;
 wire \i_ibex/ex_block_i/alu_i/_0086_ ;
 wire \i_ibex/ex_block_i/alu_i/_0087_ ;
 wire \i_ibex/ex_block_i/alu_i/_0088_ ;
 wire \i_ibex/ex_block_i/alu_i/_0089_ ;
 wire \i_ibex/ex_block_i/alu_i/_0090_ ;
 wire \i_ibex/ex_block_i/alu_i/_0091_ ;
 wire net736;
 wire \i_ibex/ex_block_i/alu_i/_0093_ ;
 wire \i_ibex/ex_block_i/alu_i/_0094_ ;
 wire net735;
 wire \i_ibex/ex_block_i/alu_i/_0096_ ;
 wire \i_ibex/ex_block_i/alu_i/_0097_ ;
 wire \i_ibex/ex_block_i/alu_i/_0098_ ;
 wire \i_ibex/ex_block_i/alu_i/_0099_ ;
 wire \i_ibex/ex_block_i/alu_i/_0100_ ;
 wire \i_ibex/ex_block_i/alu_i/_0101_ ;
 wire \i_ibex/ex_block_i/alu_i/_0102_ ;
 wire \i_ibex/ex_block_i/alu_i/_0103_ ;
 wire \i_ibex/ex_block_i/alu_i/_0104_ ;
 wire \i_ibex/ex_block_i/alu_i/_0105_ ;
 wire net734;
 wire net733;
 wire net732;
 wire net731;
 wire \i_ibex/ex_block_i/alu_i/_0110_ ;
 wire \i_ibex/ex_block_i/alu_i/_0111_ ;
 wire \i_ibex/ex_block_i/alu_i/_0112_ ;
 wire \i_ibex/ex_block_i/alu_i/_0113_ ;
 wire net730;
 wire net729;
 wire \i_ibex/ex_block_i/alu_i/_0116_ ;
 wire \i_ibex/ex_block_i/alu_i/_0117_ ;
 wire \i_ibex/ex_block_i/alu_i/_0118_ ;
 wire \i_ibex/ex_block_i/alu_i/_0119_ ;
 wire \i_ibex/ex_block_i/alu_i/_0120_ ;
 wire \i_ibex/ex_block_i/alu_i/_0121_ ;
 wire \i_ibex/ex_block_i/alu_i/_0122_ ;
 wire \i_ibex/ex_block_i/alu_i/_0123_ ;
 wire \i_ibex/ex_block_i/alu_i/_0124_ ;
 wire \i_ibex/ex_block_i/alu_i/_0125_ ;
 wire net728;
 wire \i_ibex/ex_block_i/alu_i/_0127_ ;
 wire \i_ibex/ex_block_i/alu_i/_0128_ ;
 wire \i_ibex/ex_block_i/alu_i/_0129_ ;
 wire \i_ibex/ex_block_i/alu_i/_0130_ ;
 wire \i_ibex/ex_block_i/alu_i/_0131_ ;
 wire \i_ibex/ex_block_i/alu_i/_0132_ ;
 wire \i_ibex/ex_block_i/alu_i/_0133_ ;
 wire \i_ibex/ex_block_i/alu_i/_0134_ ;
 wire \i_ibex/ex_block_i/alu_i/_0135_ ;
 wire \i_ibex/ex_block_i/alu_i/_0136_ ;
 wire \i_ibex/ex_block_i/alu_i/_0137_ ;
 wire \i_ibex/ex_block_i/alu_i/_0138_ ;
 wire \i_ibex/ex_block_i/alu_i/_0139_ ;
 wire \i_ibex/ex_block_i/alu_i/_0140_ ;
 wire \i_ibex/ex_block_i/alu_i/_0141_ ;
 wire \i_ibex/ex_block_i/alu_i/_0142_ ;
 wire \i_ibex/ex_block_i/alu_i/_0143_ ;
 wire \i_ibex/ex_block_i/alu_i/_0144_ ;
 wire \i_ibex/ex_block_i/alu_i/_0145_ ;
 wire net727;
 wire net726;
 wire \i_ibex/ex_block_i/alu_i/_0148_ ;
 wire \i_ibex/ex_block_i/alu_i/_0149_ ;
 wire \i_ibex/ex_block_i/alu_i/_0150_ ;
 wire net725;
 wire \i_ibex/ex_block_i/alu_i/_0152_ ;
 wire net724;
 wire \i_ibex/ex_block_i/alu_i/_0154_ ;
 wire net723;
 wire \i_ibex/ex_block_i/alu_i/_0156_ ;
 wire net722;
 wire \i_ibex/ex_block_i/alu_i/_0158_ ;
 wire net721;
 wire \i_ibex/ex_block_i/alu_i/_0160_ ;
 wire \i_ibex/ex_block_i/alu_i/_0161_ ;
 wire \i_ibex/ex_block_i/alu_i/_0162_ ;
 wire net720;
 wire \i_ibex/ex_block_i/alu_i/_0164_ ;
 wire net719;
 wire net718;
 wire net717;
 wire \i_ibex/ex_block_i/alu_i/_0168_ ;
 wire \i_ibex/ex_block_i/alu_i/_0169_ ;
 wire \i_ibex/ex_block_i/alu_i/_0170_ ;
 wire \i_ibex/ex_block_i/alu_i/_0171_ ;
 wire net716;
 wire net715;
 wire \i_ibex/ex_block_i/alu_i/_0174_ ;
 wire \i_ibex/ex_block_i/alu_i/_0175_ ;
 wire \i_ibex/ex_block_i/alu_i/_0176_ ;
 wire \i_ibex/ex_block_i/alu_i/_0177_ ;
 wire net714;
 wire \i_ibex/ex_block_i/alu_i/_0179_ ;
 wire net713;
 wire \i_ibex/ex_block_i/alu_i/_0181_ ;
 wire \i_ibex/ex_block_i/alu_i/_0182_ ;
 wire \i_ibex/ex_block_i/alu_i/_0183_ ;
 wire net712;
 wire \i_ibex/ex_block_i/alu_i/_0185_ ;
 wire \i_ibex/ex_block_i/alu_i/_0186_ ;
 wire \i_ibex/ex_block_i/alu_i/_0187_ ;
 wire \i_ibex/ex_block_i/alu_i/_0188_ ;
 wire \i_ibex/ex_block_i/alu_i/_0189_ ;
 wire \i_ibex/ex_block_i/alu_i/_0190_ ;
 wire \i_ibex/ex_block_i/alu_i/_0191_ ;
 wire \i_ibex/ex_block_i/alu_i/_0192_ ;
 wire \i_ibex/ex_block_i/alu_i/_0193_ ;
 wire \i_ibex/ex_block_i/alu_i/_0194_ ;
 wire \i_ibex/ex_block_i/alu_i/_0195_ ;
 wire \i_ibex/ex_block_i/alu_i/_0196_ ;
 wire \i_ibex/ex_block_i/alu_i/_0197_ ;
 wire \i_ibex/ex_block_i/alu_i/_0198_ ;
 wire \i_ibex/ex_block_i/alu_i/_0199_ ;
 wire \i_ibex/ex_block_i/alu_i/_0200_ ;
 wire \i_ibex/ex_block_i/alu_i/_0201_ ;
 wire \i_ibex/ex_block_i/alu_i/_0202_ ;
 wire \i_ibex/ex_block_i/alu_i/_0203_ ;
 wire \i_ibex/ex_block_i/alu_i/_0204_ ;
 wire \i_ibex/ex_block_i/alu_i/_0205_ ;
 wire net711;
 wire \i_ibex/ex_block_i/alu_i/_0207_ ;
 wire \i_ibex/ex_block_i/alu_i/_0208_ ;
 wire \i_ibex/ex_block_i/alu_i/_0209_ ;
 wire \i_ibex/ex_block_i/alu_i/_0210_ ;
 wire \i_ibex/ex_block_i/alu_i/_0211_ ;
 wire \i_ibex/ex_block_i/alu_i/_0212_ ;
 wire \i_ibex/ex_block_i/alu_i/_0213_ ;
 wire \i_ibex/ex_block_i/alu_i/_0214_ ;
 wire \i_ibex/ex_block_i/alu_i/_0215_ ;
 wire \i_ibex/ex_block_i/alu_i/_0216_ ;
 wire \i_ibex/ex_block_i/alu_i/_0217_ ;
 wire \i_ibex/ex_block_i/alu_i/_0218_ ;
 wire \i_ibex/ex_block_i/alu_i/_0219_ ;
 wire \i_ibex/ex_block_i/alu_i/_0220_ ;
 wire \i_ibex/ex_block_i/alu_i/_0221_ ;
 wire \i_ibex/ex_block_i/alu_i/_0222_ ;
 wire \i_ibex/ex_block_i/alu_i/_0223_ ;
 wire \i_ibex/ex_block_i/alu_i/_0224_ ;
 wire \i_ibex/ex_block_i/alu_i/_0225_ ;
 wire \i_ibex/ex_block_i/alu_i/_0226_ ;
 wire \i_ibex/ex_block_i/alu_i/_0227_ ;
 wire net710;
 wire \i_ibex/ex_block_i/alu_i/_0229_ ;
 wire \i_ibex/ex_block_i/alu_i/_0230_ ;
 wire \i_ibex/ex_block_i/alu_i/_0231_ ;
 wire \i_ibex/ex_block_i/alu_i/_0232_ ;
 wire \i_ibex/ex_block_i/alu_i/_0233_ ;
 wire \i_ibex/ex_block_i/alu_i/_0234_ ;
 wire \i_ibex/ex_block_i/alu_i/_0235_ ;
 wire \i_ibex/ex_block_i/alu_i/_0236_ ;
 wire \i_ibex/ex_block_i/alu_i/_0237_ ;
 wire \i_ibex/ex_block_i/alu_i/_0238_ ;
 wire net709;
 wire \i_ibex/ex_block_i/alu_i/_0240_ ;
 wire \i_ibex/ex_block_i/alu_i/_0241_ ;
 wire \i_ibex/ex_block_i/alu_i/_0242_ ;
 wire \i_ibex/ex_block_i/alu_i/_0243_ ;
 wire net708;
 wire \i_ibex/ex_block_i/alu_i/_0245_ ;
 wire \i_ibex/ex_block_i/alu_i/_0246_ ;
 wire \i_ibex/ex_block_i/alu_i/_0247_ ;
 wire \i_ibex/ex_block_i/alu_i/_0248_ ;
 wire \i_ibex/ex_block_i/alu_i/_0249_ ;
 wire net707;
 wire \i_ibex/ex_block_i/alu_i/_0251_ ;
 wire \i_ibex/ex_block_i/alu_i/_0252_ ;
 wire \i_ibex/ex_block_i/alu_i/_0253_ ;
 wire \i_ibex/ex_block_i/alu_i/_0254_ ;
 wire \i_ibex/ex_block_i/alu_i/_0255_ ;
 wire \i_ibex/ex_block_i/alu_i/_0256_ ;
 wire \i_ibex/ex_block_i/alu_i/_0257_ ;
 wire \i_ibex/ex_block_i/alu_i/_0258_ ;
 wire \i_ibex/ex_block_i/alu_i/_0259_ ;
 wire \i_ibex/ex_block_i/alu_i/_0260_ ;
 wire \i_ibex/ex_block_i/alu_i/_0261_ ;
 wire \i_ibex/ex_block_i/alu_i/_0262_ ;
 wire \i_ibex/ex_block_i/alu_i/_0263_ ;
 wire \i_ibex/ex_block_i/alu_i/_0264_ ;
 wire \i_ibex/ex_block_i/alu_i/_0265_ ;
 wire \i_ibex/ex_block_i/alu_i/_0266_ ;
 wire \i_ibex/ex_block_i/alu_i/_0267_ ;
 wire \i_ibex/ex_block_i/alu_i/_0268_ ;
 wire \i_ibex/ex_block_i/alu_i/_0269_ ;
 wire \i_ibex/ex_block_i/alu_i/_0270_ ;
 wire \i_ibex/ex_block_i/alu_i/_0271_ ;
 wire \i_ibex/ex_block_i/alu_i/_0272_ ;
 wire \i_ibex/ex_block_i/alu_i/_0273_ ;
 wire \i_ibex/ex_block_i/alu_i/_0274_ ;
 wire \i_ibex/ex_block_i/alu_i/_0275_ ;
 wire \i_ibex/ex_block_i/alu_i/_0276_ ;
 wire \i_ibex/ex_block_i/alu_i/_0277_ ;
 wire \i_ibex/ex_block_i/alu_i/_0278_ ;
 wire \i_ibex/ex_block_i/alu_i/_0279_ ;
 wire \i_ibex/ex_block_i/alu_i/_0280_ ;
 wire \i_ibex/ex_block_i/alu_i/_0281_ ;
 wire \i_ibex/ex_block_i/alu_i/_0282_ ;
 wire \i_ibex/ex_block_i/alu_i/_0283_ ;
 wire \i_ibex/ex_block_i/alu_i/_0284_ ;
 wire \i_ibex/ex_block_i/alu_i/_0285_ ;
 wire \i_ibex/ex_block_i/alu_i/_0286_ ;
 wire \i_ibex/ex_block_i/alu_i/_0287_ ;
 wire \i_ibex/ex_block_i/alu_i/_0288_ ;
 wire \i_ibex/ex_block_i/alu_i/_0289_ ;
 wire \i_ibex/ex_block_i/alu_i/_0290_ ;
 wire \i_ibex/ex_block_i/alu_i/_0291_ ;
 wire \i_ibex/ex_block_i/alu_i/_0292_ ;
 wire \i_ibex/ex_block_i/alu_i/_0293_ ;
 wire \i_ibex/ex_block_i/alu_i/_0294_ ;
 wire \i_ibex/ex_block_i/alu_i/_0295_ ;
 wire \i_ibex/ex_block_i/alu_i/_0296_ ;
 wire \i_ibex/ex_block_i/alu_i/_0297_ ;
 wire \i_ibex/ex_block_i/alu_i/_0298_ ;
 wire \i_ibex/ex_block_i/alu_i/_0299_ ;
 wire \i_ibex/ex_block_i/alu_i/_0300_ ;
 wire \i_ibex/ex_block_i/alu_i/_0301_ ;
 wire \i_ibex/ex_block_i/alu_i/_0302_ ;
 wire \i_ibex/ex_block_i/alu_i/_0303_ ;
 wire \i_ibex/ex_block_i/alu_i/_0304_ ;
 wire \i_ibex/ex_block_i/alu_i/_0305_ ;
 wire \i_ibex/ex_block_i/alu_i/_0306_ ;
 wire \i_ibex/ex_block_i/alu_i/_0307_ ;
 wire \i_ibex/ex_block_i/alu_i/_0308_ ;
 wire \i_ibex/ex_block_i/alu_i/_0309_ ;
 wire \i_ibex/ex_block_i/alu_i/_0310_ ;
 wire \i_ibex/ex_block_i/alu_i/_0311_ ;
 wire \i_ibex/ex_block_i/alu_i/_0312_ ;
 wire \i_ibex/ex_block_i/alu_i/_0313_ ;
 wire \i_ibex/ex_block_i/alu_i/_0314_ ;
 wire \i_ibex/ex_block_i/alu_i/_0315_ ;
 wire \i_ibex/ex_block_i/alu_i/_0316_ ;
 wire \i_ibex/ex_block_i/alu_i/_0317_ ;
 wire \i_ibex/ex_block_i/alu_i/_0318_ ;
 wire \i_ibex/ex_block_i/alu_i/_0319_ ;
 wire \i_ibex/ex_block_i/alu_i/_0320_ ;
 wire \i_ibex/ex_block_i/alu_i/_0321_ ;
 wire \i_ibex/ex_block_i/alu_i/_0322_ ;
 wire \i_ibex/ex_block_i/alu_i/_0323_ ;
 wire \i_ibex/ex_block_i/alu_i/_0324_ ;
 wire \i_ibex/ex_block_i/alu_i/_0325_ ;
 wire \i_ibex/ex_block_i/alu_i/_0326_ ;
 wire \i_ibex/ex_block_i/alu_i/_0327_ ;
 wire \i_ibex/ex_block_i/alu_i/_0328_ ;
 wire \i_ibex/ex_block_i/alu_i/_0329_ ;
 wire \i_ibex/ex_block_i/alu_i/_0330_ ;
 wire \i_ibex/ex_block_i/alu_i/_0331_ ;
 wire \i_ibex/ex_block_i/alu_i/_0332_ ;
 wire \i_ibex/ex_block_i/alu_i/_0333_ ;
 wire net706;
 wire net705;
 wire \i_ibex/ex_block_i/alu_i/_0336_ ;
 wire \i_ibex/ex_block_i/alu_i/_0337_ ;
 wire \i_ibex/ex_block_i/alu_i/_0338_ ;
 wire \i_ibex/ex_block_i/alu_i/_0339_ ;
 wire \i_ibex/ex_block_i/alu_i/_0340_ ;
 wire net704;
 wire \i_ibex/ex_block_i/alu_i/_0342_ ;
 wire net703;
 wire \i_ibex/ex_block_i/alu_i/_0344_ ;
 wire \i_ibex/ex_block_i/alu_i/_0345_ ;
 wire \i_ibex/ex_block_i/alu_i/_0346_ ;
 wire \i_ibex/ex_block_i/alu_i/_0347_ ;
 wire \i_ibex/ex_block_i/alu_i/_0348_ ;
 wire \i_ibex/ex_block_i/alu_i/_0349_ ;
 wire net702;
 wire net701;
 wire net700;
 wire \i_ibex/ex_block_i/alu_i/_0353_ ;
 wire \i_ibex/ex_block_i/alu_i/_0354_ ;
 wire \i_ibex/ex_block_i/alu_i/_0355_ ;
 wire \i_ibex/ex_block_i/alu_i/_0356_ ;
 wire \i_ibex/ex_block_i/alu_i/_0357_ ;
 wire net699;
 wire \i_ibex/ex_block_i/alu_i/_0359_ ;
 wire \i_ibex/ex_block_i/alu_i/_0360_ ;
 wire \i_ibex/ex_block_i/alu_i/_0361_ ;
 wire \i_ibex/ex_block_i/alu_i/_0362_ ;
 wire net698;
 wire \i_ibex/ex_block_i/alu_i/_0364_ ;
 wire net697;
 wire \i_ibex/ex_block_i/alu_i/_0366_ ;
 wire \i_ibex/ex_block_i/alu_i/_0367_ ;
 wire \i_ibex/ex_block_i/alu_i/_0368_ ;
 wire \i_ibex/ex_block_i/alu_i/_0369_ ;
 wire \i_ibex/ex_block_i/alu_i/_0370_ ;
 wire \i_ibex/ex_block_i/alu_i/_0371_ ;
 wire \i_ibex/ex_block_i/alu_i/_0372_ ;
 wire \i_ibex/ex_block_i/alu_i/_0373_ ;
 wire \i_ibex/ex_block_i/alu_i/_0374_ ;
 wire \i_ibex/ex_block_i/alu_i/_0375_ ;
 wire \i_ibex/ex_block_i/alu_i/_0376_ ;
 wire \i_ibex/ex_block_i/alu_i/_0377_ ;
 wire \i_ibex/ex_block_i/alu_i/_0378_ ;
 wire \i_ibex/ex_block_i/alu_i/_0379_ ;
 wire \i_ibex/ex_block_i/alu_i/_0380_ ;
 wire \i_ibex/ex_block_i/alu_i/_0381_ ;
 wire \i_ibex/ex_block_i/alu_i/_0382_ ;
 wire \i_ibex/ex_block_i/alu_i/_0383_ ;
 wire \i_ibex/ex_block_i/alu_i/_0384_ ;
 wire \i_ibex/ex_block_i/alu_i/_0385_ ;
 wire \i_ibex/ex_block_i/alu_i/_0386_ ;
 wire net696;
 wire \i_ibex/ex_block_i/alu_i/_0388_ ;
 wire \i_ibex/ex_block_i/alu_i/_0389_ ;
 wire \i_ibex/ex_block_i/alu_i/_0390_ ;
 wire \i_ibex/ex_block_i/alu_i/_0391_ ;
 wire \i_ibex/ex_block_i/alu_i/_0392_ ;
 wire \i_ibex/ex_block_i/alu_i/_0393_ ;
 wire \i_ibex/ex_block_i/alu_i/_0394_ ;
 wire \i_ibex/ex_block_i/alu_i/_0395_ ;
 wire \i_ibex/ex_block_i/alu_i/_0396_ ;
 wire \i_ibex/ex_block_i/alu_i/_0397_ ;
 wire \i_ibex/ex_block_i/alu_i/_0398_ ;
 wire \i_ibex/ex_block_i/alu_i/_0399_ ;
 wire \i_ibex/ex_block_i/alu_i/_0400_ ;
 wire \i_ibex/ex_block_i/alu_i/_0401_ ;
 wire \i_ibex/ex_block_i/alu_i/_0402_ ;
 wire \i_ibex/ex_block_i/alu_i/_0403_ ;
 wire \i_ibex/ex_block_i/alu_i/_0404_ ;
 wire \i_ibex/ex_block_i/alu_i/_0405_ ;
 wire \i_ibex/ex_block_i/alu_i/_0406_ ;
 wire \i_ibex/ex_block_i/alu_i/_0407_ ;
 wire \i_ibex/ex_block_i/alu_i/_0408_ ;
 wire \i_ibex/ex_block_i/alu_i/_0409_ ;
 wire \i_ibex/ex_block_i/alu_i/_0410_ ;
 wire \i_ibex/ex_block_i/alu_i/_0411_ ;
 wire \i_ibex/ex_block_i/alu_i/_0412_ ;
 wire \i_ibex/ex_block_i/alu_i/_0413_ ;
 wire \i_ibex/ex_block_i/alu_i/_0414_ ;
 wire \i_ibex/ex_block_i/alu_i/_0415_ ;
 wire \i_ibex/ex_block_i/alu_i/_0416_ ;
 wire \i_ibex/ex_block_i/alu_i/_0417_ ;
 wire \i_ibex/ex_block_i/alu_i/_0418_ ;
 wire \i_ibex/ex_block_i/alu_i/_0419_ ;
 wire \i_ibex/ex_block_i/alu_i/_0420_ ;
 wire \i_ibex/ex_block_i/alu_i/_0421_ ;
 wire \i_ibex/ex_block_i/alu_i/_0422_ ;
 wire \i_ibex/ex_block_i/alu_i/_0423_ ;
 wire \i_ibex/ex_block_i/alu_i/_0424_ ;
 wire \i_ibex/ex_block_i/alu_i/_0425_ ;
 wire \i_ibex/ex_block_i/alu_i/_0426_ ;
 wire \i_ibex/ex_block_i/alu_i/_0427_ ;
 wire \i_ibex/ex_block_i/alu_i/_0428_ ;
 wire \i_ibex/ex_block_i/alu_i/_0429_ ;
 wire \i_ibex/ex_block_i/alu_i/_0430_ ;
 wire \i_ibex/ex_block_i/alu_i/_0431_ ;
 wire \i_ibex/ex_block_i/alu_i/_0432_ ;
 wire \i_ibex/ex_block_i/alu_i/_0433_ ;
 wire \i_ibex/ex_block_i/alu_i/_0434_ ;
 wire \i_ibex/ex_block_i/alu_i/_0435_ ;
 wire \i_ibex/ex_block_i/alu_i/_0436_ ;
 wire \i_ibex/ex_block_i/alu_i/_0437_ ;
 wire \i_ibex/ex_block_i/alu_i/_0438_ ;
 wire \i_ibex/ex_block_i/alu_i/_0439_ ;
 wire \i_ibex/ex_block_i/alu_i/_0440_ ;
 wire \i_ibex/ex_block_i/alu_i/_0441_ ;
 wire \i_ibex/ex_block_i/alu_i/_0442_ ;
 wire \i_ibex/ex_block_i/alu_i/_0443_ ;
 wire \i_ibex/ex_block_i/alu_i/_0444_ ;
 wire \i_ibex/ex_block_i/alu_i/_0445_ ;
 wire \i_ibex/ex_block_i/alu_i/_0446_ ;
 wire \i_ibex/ex_block_i/alu_i/_0447_ ;
 wire \i_ibex/ex_block_i/alu_i/_0448_ ;
 wire \i_ibex/ex_block_i/alu_i/_0449_ ;
 wire \i_ibex/ex_block_i/alu_i/_0450_ ;
 wire \i_ibex/ex_block_i/alu_i/_0451_ ;
 wire \i_ibex/ex_block_i/alu_i/_0452_ ;
 wire \i_ibex/ex_block_i/alu_i/_0453_ ;
 wire \i_ibex/ex_block_i/alu_i/_0454_ ;
 wire \i_ibex/ex_block_i/alu_i/_0455_ ;
 wire \i_ibex/ex_block_i/alu_i/_0456_ ;
 wire \i_ibex/ex_block_i/alu_i/_0457_ ;
 wire \i_ibex/ex_block_i/alu_i/_0458_ ;
 wire \i_ibex/ex_block_i/alu_i/_0459_ ;
 wire \i_ibex/ex_block_i/alu_i/_0460_ ;
 wire \i_ibex/ex_block_i/alu_i/_0461_ ;
 wire \i_ibex/ex_block_i/alu_i/_0462_ ;
 wire \i_ibex/ex_block_i/alu_i/_0463_ ;
 wire \i_ibex/ex_block_i/alu_i/_0464_ ;
 wire \i_ibex/ex_block_i/alu_i/_0465_ ;
 wire \i_ibex/ex_block_i/alu_i/_0466_ ;
 wire \i_ibex/ex_block_i/alu_i/_0467_ ;
 wire \i_ibex/ex_block_i/alu_i/_0468_ ;
 wire \i_ibex/ex_block_i/alu_i/_0469_ ;
 wire net695;
 wire net694;
 wire net693;
 wire \i_ibex/ex_block_i/alu_i/_0473_ ;
 wire \i_ibex/ex_block_i/alu_i/_0474_ ;
 wire \i_ibex/ex_block_i/alu_i/_0475_ ;
 wire \i_ibex/ex_block_i/alu_i/_0476_ ;
 wire \i_ibex/ex_block_i/alu_i/_0477_ ;
 wire \i_ibex/ex_block_i/alu_i/_0478_ ;
 wire \i_ibex/ex_block_i/alu_i/_0479_ ;
 wire \i_ibex/ex_block_i/alu_i/_0480_ ;
 wire \i_ibex/ex_block_i/alu_i/_0481_ ;
 wire \i_ibex/ex_block_i/alu_i/_0482_ ;
 wire net692;
 wire \i_ibex/ex_block_i/alu_i/_0484_ ;
 wire \i_ibex/ex_block_i/alu_i/_0485_ ;
 wire \i_ibex/ex_block_i/alu_i/_0486_ ;
 wire \i_ibex/ex_block_i/alu_i/_0487_ ;
 wire \i_ibex/ex_block_i/alu_i/_0488_ ;
 wire \i_ibex/ex_block_i/alu_i/_0489_ ;
 wire \i_ibex/ex_block_i/alu_i/_0490_ ;
 wire \i_ibex/ex_block_i/alu_i/_0491_ ;
 wire \i_ibex/ex_block_i/alu_i/_0492_ ;
 wire \i_ibex/ex_block_i/alu_i/_0493_ ;
 wire \i_ibex/ex_block_i/alu_i/_0494_ ;
 wire \i_ibex/ex_block_i/alu_i/_0495_ ;
 wire \i_ibex/ex_block_i/alu_i/_0496_ ;
 wire \i_ibex/ex_block_i/alu_i/_0497_ ;
 wire \i_ibex/ex_block_i/alu_i/_0498_ ;
 wire \i_ibex/ex_block_i/alu_i/_0499_ ;
 wire \i_ibex/ex_block_i/alu_i/_0500_ ;
 wire \i_ibex/ex_block_i/alu_i/_0501_ ;
 wire \i_ibex/ex_block_i/alu_i/_0502_ ;
 wire \i_ibex/ex_block_i/alu_i/_0503_ ;
 wire \i_ibex/ex_block_i/alu_i/_0504_ ;
 wire \i_ibex/ex_block_i/alu_i/_0505_ ;
 wire \i_ibex/ex_block_i/alu_i/_0506_ ;
 wire \i_ibex/ex_block_i/alu_i/_0507_ ;
 wire \i_ibex/ex_block_i/alu_i/_0508_ ;
 wire \i_ibex/ex_block_i/alu_i/_0509_ ;
 wire \i_ibex/ex_block_i/alu_i/_0510_ ;
 wire \i_ibex/ex_block_i/alu_i/_0511_ ;
 wire \i_ibex/ex_block_i/alu_i/_0512_ ;
 wire \i_ibex/ex_block_i/alu_i/_0513_ ;
 wire \i_ibex/ex_block_i/alu_i/_0514_ ;
 wire \i_ibex/ex_block_i/alu_i/_0515_ ;
 wire \i_ibex/ex_block_i/alu_i/_0516_ ;
 wire \i_ibex/ex_block_i/alu_i/_0517_ ;
 wire \i_ibex/ex_block_i/alu_i/_0518_ ;
 wire \i_ibex/ex_block_i/alu_i/_0519_ ;
 wire \i_ibex/ex_block_i/alu_i/_0520_ ;
 wire \i_ibex/ex_block_i/alu_i/_0521_ ;
 wire \i_ibex/ex_block_i/alu_i/_0522_ ;
 wire \i_ibex/ex_block_i/alu_i/_0523_ ;
 wire \i_ibex/ex_block_i/alu_i/_0524_ ;
 wire \i_ibex/ex_block_i/alu_i/_0525_ ;
 wire \i_ibex/ex_block_i/alu_i/_0526_ ;
 wire \i_ibex/ex_block_i/alu_i/_0527_ ;
 wire \i_ibex/ex_block_i/alu_i/_0528_ ;
 wire \i_ibex/ex_block_i/alu_i/_0529_ ;
 wire \i_ibex/ex_block_i/alu_i/_0530_ ;
 wire \i_ibex/ex_block_i/alu_i/_0531_ ;
 wire \i_ibex/ex_block_i/alu_i/_0532_ ;
 wire \i_ibex/ex_block_i/alu_i/_0533_ ;
 wire \i_ibex/ex_block_i/alu_i/_0534_ ;
 wire \i_ibex/ex_block_i/alu_i/_0535_ ;
 wire \i_ibex/ex_block_i/alu_i/_0536_ ;
 wire \i_ibex/ex_block_i/alu_i/_0537_ ;
 wire \i_ibex/ex_block_i/alu_i/_0538_ ;
 wire \i_ibex/ex_block_i/alu_i/_0539_ ;
 wire \i_ibex/ex_block_i/alu_i/_0540_ ;
 wire \i_ibex/ex_block_i/alu_i/_0541_ ;
 wire \i_ibex/ex_block_i/alu_i/_0542_ ;
 wire \i_ibex/ex_block_i/alu_i/_0543_ ;
 wire \i_ibex/ex_block_i/alu_i/_0544_ ;
 wire \i_ibex/ex_block_i/alu_i/_0545_ ;
 wire \i_ibex/ex_block_i/alu_i/_0546_ ;
 wire \i_ibex/ex_block_i/alu_i/_0547_ ;
 wire \i_ibex/ex_block_i/alu_i/_0548_ ;
 wire \i_ibex/ex_block_i/alu_i/_0549_ ;
 wire \i_ibex/ex_block_i/alu_i/_0550_ ;
 wire \i_ibex/ex_block_i/alu_i/_0551_ ;
 wire \i_ibex/ex_block_i/alu_i/_0552_ ;
 wire \i_ibex/ex_block_i/alu_i/_0553_ ;
 wire \i_ibex/ex_block_i/alu_i/_0554_ ;
 wire \i_ibex/ex_block_i/alu_i/_0555_ ;
 wire \i_ibex/ex_block_i/alu_i/_0556_ ;
 wire \i_ibex/ex_block_i/alu_i/_0557_ ;
 wire \i_ibex/ex_block_i/alu_i/_0558_ ;
 wire \i_ibex/ex_block_i/alu_i/_0559_ ;
 wire \i_ibex/ex_block_i/alu_i/_0560_ ;
 wire \i_ibex/ex_block_i/alu_i/_0561_ ;
 wire \i_ibex/ex_block_i/alu_i/_0562_ ;
 wire \i_ibex/ex_block_i/alu_i/_0563_ ;
 wire \i_ibex/ex_block_i/alu_i/_0564_ ;
 wire \i_ibex/ex_block_i/alu_i/_0565_ ;
 wire \i_ibex/ex_block_i/alu_i/_0566_ ;
 wire \i_ibex/ex_block_i/alu_i/_0567_ ;
 wire \i_ibex/ex_block_i/alu_i/_0568_ ;
 wire \i_ibex/ex_block_i/alu_i/_0569_ ;
 wire \i_ibex/ex_block_i/alu_i/_0570_ ;
 wire \i_ibex/ex_block_i/alu_i/_0571_ ;
 wire \i_ibex/ex_block_i/alu_i/_0572_ ;
 wire \i_ibex/ex_block_i/alu_i/_0573_ ;
 wire \i_ibex/ex_block_i/alu_i/_0574_ ;
 wire \i_ibex/ex_block_i/alu_i/_0575_ ;
 wire \i_ibex/ex_block_i/alu_i/_0576_ ;
 wire \i_ibex/ex_block_i/alu_i/_0577_ ;
 wire \i_ibex/ex_block_i/alu_i/_0578_ ;
 wire \i_ibex/ex_block_i/alu_i/_0579_ ;
 wire \i_ibex/ex_block_i/alu_i/_0580_ ;
 wire \i_ibex/ex_block_i/alu_i/_0581_ ;
 wire \i_ibex/ex_block_i/alu_i/_0582_ ;
 wire \i_ibex/ex_block_i/alu_i/_0583_ ;
 wire \i_ibex/ex_block_i/alu_i/_0584_ ;
 wire \i_ibex/ex_block_i/alu_i/_0585_ ;
 wire \i_ibex/ex_block_i/alu_i/_0586_ ;
 wire \i_ibex/ex_block_i/alu_i/_0587_ ;
 wire \i_ibex/ex_block_i/alu_i/_0588_ ;
 wire \i_ibex/ex_block_i/alu_i/_0589_ ;
 wire net826;
 wire net825;
 wire net824;
 wire net823;
 wire net822;
 wire net821;
 wire net820;
 wire \i_ibex/ex_block_i/alu_i/_0597_ ;
 wire net819;
 wire net818;
 wire \i_ibex/ex_block_i/alu_i/_0600_ ;
 wire \i_ibex/ex_block_i/alu_i/_0601_ ;
 wire net817;
 wire \i_ibex/ex_block_i/alu_i/_0603_ ;
 wire \i_ibex/ex_block_i/alu_i/_0604_ ;
 wire \i_ibex/ex_block_i/alu_i/_0605_ ;
 wire \i_ibex/ex_block_i/alu_i/_0606_ ;
 wire \i_ibex/ex_block_i/alu_i/_0607_ ;
 wire \i_ibex/ex_block_i/alu_i/_0608_ ;
 wire net816;
 wire \i_ibex/ex_block_i/alu_i/_0610_ ;
 wire \i_ibex/ex_block_i/alu_i/_0611_ ;
 wire \i_ibex/ex_block_i/alu_i/_0612_ ;
 wire net815;
 wire \i_ibex/ex_block_i/alu_i/_0614_ ;
 wire \i_ibex/ex_block_i/alu_i/_0615_ ;
 wire \i_ibex/ex_block_i/alu_i/_0616_ ;
 wire \i_ibex/ex_block_i/alu_i/_0617_ ;
 wire \i_ibex/ex_block_i/alu_i/_0618_ ;
 wire \i_ibex/ex_block_i/alu_i/_0619_ ;
 wire \i_ibex/ex_block_i/alu_i/_0620_ ;
 wire \i_ibex/ex_block_i/alu_i/_0621_ ;
 wire net814;
 wire net813;
 wire net812;
 wire net811;
 wire \i_ibex/ex_block_i/alu_i/_0626_ ;
 wire \i_ibex/ex_block_i/alu_i/_0627_ ;
 wire net810;
 wire net809;
 wire net808;
 wire net807;
 wire net806;
 wire net805;
 wire net804;
 wire \i_ibex/ex_block_i/alu_i/_0635_ ;
 wire \i_ibex/ex_block_i/alu_i/_0636_ ;
 wire \i_ibex/ex_block_i/alu_i/_0637_ ;
 wire \i_ibex/ex_block_i/alu_i/_0638_ ;
 wire \i_ibex/ex_block_i/alu_i/_0639_ ;
 wire net803;
 wire \i_ibex/ex_block_i/alu_i/_0641_ ;
 wire \i_ibex/ex_block_i/alu_i/_0642_ ;
 wire \i_ibex/ex_block_i/alu_i/_0643_ ;
 wire \i_ibex/ex_block_i/alu_i/_0644_ ;
 wire \i_ibex/ex_block_i/alu_i/_0645_ ;
 wire \i_ibex/ex_block_i/alu_i/_0646_ ;
 wire \i_ibex/ex_block_i/alu_i/_0647_ ;
 wire \i_ibex/ex_block_i/alu_i/_0648_ ;
 wire \i_ibex/ex_block_i/alu_i/_0649_ ;
 wire \i_ibex/ex_block_i/alu_i/_0650_ ;
 wire net802;
 wire \i_ibex/ex_block_i/alu_i/_0652_ ;
 wire \i_ibex/ex_block_i/alu_i/_0653_ ;
 wire \i_ibex/ex_block_i/alu_i/_0654_ ;
 wire \i_ibex/ex_block_i/alu_i/_0655_ ;
 wire \i_ibex/ex_block_i/alu_i/_0656_ ;
 wire \i_ibex/ex_block_i/alu_i/_0657_ ;
 wire \i_ibex/ex_block_i/alu_i/_0658_ ;
 wire net801;
 wire \i_ibex/ex_block_i/alu_i/_0660_ ;
 wire \i_ibex/ex_block_i/alu_i/_0661_ ;
 wire \i_ibex/ex_block_i/alu_i/_0662_ ;
 wire \i_ibex/ex_block_i/alu_i/_0663_ ;
 wire \i_ibex/ex_block_i/alu_i/_0664_ ;
 wire \i_ibex/ex_block_i/alu_i/_0665_ ;
 wire net800;
 wire \i_ibex/ex_block_i/alu_i/_0667_ ;
 wire \i_ibex/ex_block_i/alu_i/_0668_ ;
 wire \i_ibex/ex_block_i/alu_i/_0669_ ;
 wire \i_ibex/ex_block_i/alu_i/_0670_ ;
 wire \i_ibex/ex_block_i/alu_i/_0671_ ;
 wire \i_ibex/ex_block_i/alu_i/_0672_ ;
 wire net799;
 wire \i_ibex/ex_block_i/alu_i/_0674_ ;
 wire \i_ibex/ex_block_i/alu_i/_0675_ ;
 wire \i_ibex/ex_block_i/alu_i/_0676_ ;
 wire \i_ibex/ex_block_i/alu_i/_0677_ ;
 wire net798;
 wire net797;
 wire \i_ibex/ex_block_i/alu_i/_0680_ ;
 wire \i_ibex/ex_block_i/alu_i/_0681_ ;
 wire \i_ibex/ex_block_i/alu_i/_0682_ ;
 wire net796;
 wire \i_ibex/ex_block_i/alu_i/_0684_ ;
 wire \i_ibex/ex_block_i/alu_i/_0685_ ;
 wire \i_ibex/ex_block_i/alu_i/_0686_ ;
 wire \i_ibex/ex_block_i/alu_i/_0687_ ;
 wire \i_ibex/ex_block_i/alu_i/_0688_ ;
 wire \i_ibex/ex_block_i/alu_i/_0689_ ;
 wire \i_ibex/ex_block_i/alu_i/_0690_ ;
 wire net795;
 wire \i_ibex/ex_block_i/alu_i/_0692_ ;
 wire \i_ibex/ex_block_i/alu_i/_0693_ ;
 wire \i_ibex/ex_block_i/alu_i/_0694_ ;
 wire \i_ibex/ex_block_i/alu_i/_0695_ ;
 wire net794;
 wire \i_ibex/ex_block_i/alu_i/_0697_ ;
 wire \i_ibex/ex_block_i/alu_i/_0698_ ;
 wire \i_ibex/ex_block_i/alu_i/_0699_ ;
 wire net793;
 wire \i_ibex/ex_block_i/alu_i/_0701_ ;
 wire \i_ibex/ex_block_i/alu_i/_0702_ ;
 wire \i_ibex/ex_block_i/alu_i/_0703_ ;
 wire \i_ibex/ex_block_i/alu_i/_0704_ ;
 wire \i_ibex/ex_block_i/alu_i/_0705_ ;
 wire \i_ibex/ex_block_i/alu_i/_0706_ ;
 wire net792;
 wire net791;
 wire net790;
 wire net789;
 wire \i_ibex/ex_block_i/alu_i/_0711_ ;
 wire \i_ibex/ex_block_i/alu_i/_0712_ ;
 wire \i_ibex/ex_block_i/alu_i/_0713_ ;
 wire \i_ibex/ex_block_i/alu_i/_0714_ ;
 wire \i_ibex/ex_block_i/alu_i/_0715_ ;
 wire \i_ibex/ex_block_i/alu_i/_0716_ ;
 wire \i_ibex/ex_block_i/alu_i/_0717_ ;
 wire \i_ibex/ex_block_i/alu_i/_0718_ ;
 wire net788;
 wire \i_ibex/ex_block_i/alu_i/_0720_ ;
 wire \i_ibex/ex_block_i/alu_i/_0721_ ;
 wire net787;
 wire net786;
 wire \i_ibex/ex_block_i/alu_i/_0724_ ;
 wire \i_ibex/ex_block_i/alu_i/_0725_ ;
 wire \i_ibex/ex_block_i/alu_i/_0726_ ;
 wire \i_ibex/ex_block_i/alu_i/_0727_ ;
 wire net785;
 wire \i_ibex/ex_block_i/alu_i/_0729_ ;
 wire net784;
 wire \i_ibex/ex_block_i/alu_i/_0731_ ;
 wire \i_ibex/ex_block_i/alu_i/_0732_ ;
 wire \i_ibex/ex_block_i/alu_i/_0733_ ;
 wire \i_ibex/ex_block_i/alu_i/_0734_ ;
 wire \i_ibex/ex_block_i/alu_i/_0735_ ;
 wire \i_ibex/ex_block_i/alu_i/_0736_ ;
 wire \i_ibex/ex_block_i/alu_i/_0737_ ;
 wire \i_ibex/ex_block_i/alu_i/_0738_ ;
 wire net783;
 wire \i_ibex/ex_block_i/alu_i/_0740_ ;
 wire \i_ibex/ex_block_i/alu_i/_0741_ ;
 wire \i_ibex/ex_block_i/alu_i/_0742_ ;
 wire \i_ibex/ex_block_i/alu_i/_0743_ ;
 wire \i_ibex/ex_block_i/alu_i/_0744_ ;
 wire \i_ibex/ex_block_i/alu_i/_0745_ ;
 wire \i_ibex/ex_block_i/alu_i/_0746_ ;
 wire \i_ibex/ex_block_i/alu_i/_0747_ ;
 wire \i_ibex/ex_block_i/alu_i/_0748_ ;
 wire \i_ibex/ex_block_i/alu_i/_0749_ ;
 wire \i_ibex/ex_block_i/alu_i/_0750_ ;
 wire \i_ibex/ex_block_i/alu_i/_0751_ ;
 wire \i_ibex/ex_block_i/alu_i/_0752_ ;
 wire \i_ibex/ex_block_i/alu_i/_0753_ ;
 wire \i_ibex/ex_block_i/alu_i/_0754_ ;
 wire \i_ibex/ex_block_i/alu_i/_0755_ ;
 wire \i_ibex/ex_block_i/alu_i/_0756_ ;
 wire \i_ibex/ex_block_i/alu_i/_0757_ ;
 wire \i_ibex/ex_block_i/alu_i/_0758_ ;
 wire net782;
 wire \i_ibex/ex_block_i/alu_i/_0760_ ;
 wire net781;
 wire \i_ibex/ex_block_i/alu_i/_0762_ ;
 wire \i_ibex/ex_block_i/alu_i/_0763_ ;
 wire \i_ibex/ex_block_i/alu_i/_0764_ ;
 wire \i_ibex/ex_block_i/alu_i/_0765_ ;
 wire \i_ibex/ex_block_i/alu_i/_0766_ ;
 wire \i_ibex/ex_block_i/alu_i/_0767_ ;
 wire \i_ibex/ex_block_i/alu_i/_0768_ ;
 wire net780;
 wire net779;
 wire \i_ibex/ex_block_i/alu_i/_0771_ ;
 wire \i_ibex/ex_block_i/alu_i/_0772_ ;
 wire \i_ibex/ex_block_i/alu_i/_0773_ ;
 wire \i_ibex/ex_block_i/alu_i/_0774_ ;
 wire \i_ibex/ex_block_i/alu_i/_0775_ ;
 wire net778;
 wire \i_ibex/ex_block_i/alu_i/_0777_ ;
 wire net777;
 wire \i_ibex/ex_block_i/alu_i/_0779_ ;
 wire \i_ibex/ex_block_i/alu_i/_0780_ ;
 wire \i_ibex/ex_block_i/alu_i/_0781_ ;
 wire \i_ibex/ex_block_i/alu_i/_0782_ ;
 wire \i_ibex/ex_block_i/alu_i/_0783_ ;
 wire \i_ibex/ex_block_i/alu_i/_0784_ ;
 wire \i_ibex/ex_block_i/alu_i/_0785_ ;
 wire \i_ibex/ex_block_i/alu_i/_0786_ ;
 wire \i_ibex/ex_block_i/alu_i/_0787_ ;
 wire \i_ibex/ex_block_i/alu_i/_0788_ ;
 wire net776;
 wire \i_ibex/ex_block_i/alu_i/_0790_ ;
 wire \i_ibex/ex_block_i/alu_i/_0791_ ;
 wire net775;
 wire \i_ibex/ex_block_i/alu_i/_0793_ ;
 wire \i_ibex/ex_block_i/alu_i/_0794_ ;
 wire \i_ibex/ex_block_i/alu_i/_0795_ ;
 wire net774;
 wire net773;
 wire \i_ibex/ex_block_i/alu_i/_0798_ ;
 wire \i_ibex/ex_block_i/alu_i/_0799_ ;
 wire \i_ibex/ex_block_i/alu_i/_0800_ ;
 wire \i_ibex/ex_block_i/alu_i/_0801_ ;
 wire \i_ibex/ex_block_i/alu_i/_0802_ ;
 wire \i_ibex/ex_block_i/alu_i/_0803_ ;
 wire \i_ibex/ex_block_i/alu_i/_0804_ ;
 wire \i_ibex/ex_block_i/alu_i/_0805_ ;
 wire \i_ibex/ex_block_i/alu_i/_0806_ ;
 wire \i_ibex/ex_block_i/alu_i/_0807_ ;
 wire \i_ibex/ex_block_i/alu_i/_0808_ ;
 wire \i_ibex/ex_block_i/alu_i/_0809_ ;
 wire \i_ibex/ex_block_i/alu_i/_0810_ ;
 wire \i_ibex/ex_block_i/alu_i/_0811_ ;
 wire \i_ibex/ex_block_i/alu_i/_0812_ ;
 wire \i_ibex/ex_block_i/alu_i/_0813_ ;
 wire \i_ibex/ex_block_i/alu_i/_0814_ ;
 wire \i_ibex/ex_block_i/alu_i/_0815_ ;
 wire \i_ibex/ex_block_i/alu_i/_0816_ ;
 wire \i_ibex/ex_block_i/alu_i/_0817_ ;
 wire \i_ibex/ex_block_i/alu_i/_0818_ ;
 wire \i_ibex/ex_block_i/alu_i/_0819_ ;
 wire \i_ibex/ex_block_i/alu_i/_0820_ ;
 wire \i_ibex/ex_block_i/alu_i/_0821_ ;
 wire \i_ibex/ex_block_i/alu_i/_0822_ ;
 wire \i_ibex/ex_block_i/alu_i/_0823_ ;
 wire \i_ibex/ex_block_i/alu_i/_0824_ ;
 wire \i_ibex/ex_block_i/alu_i/_0825_ ;
 wire \i_ibex/ex_block_i/alu_i/_0826_ ;
 wire \i_ibex/ex_block_i/alu_i/_0827_ ;
 wire \i_ibex/ex_block_i/alu_i/_0828_ ;
 wire \i_ibex/ex_block_i/alu_i/_0829_ ;
 wire \i_ibex/ex_block_i/alu_i/_0830_ ;
 wire \i_ibex/ex_block_i/alu_i/_0831_ ;
 wire \i_ibex/ex_block_i/alu_i/_0832_ ;
 wire \i_ibex/ex_block_i/alu_i/_0833_ ;
 wire \i_ibex/ex_block_i/alu_i/_0834_ ;
 wire \i_ibex/ex_block_i/alu_i/_0835_ ;
 wire \i_ibex/ex_block_i/alu_i/_0836_ ;
 wire \i_ibex/ex_block_i/alu_i/_0837_ ;
 wire \i_ibex/ex_block_i/alu_i/_0838_ ;
 wire \i_ibex/ex_block_i/alu_i/_0839_ ;
 wire \i_ibex/ex_block_i/alu_i/_0840_ ;
 wire \i_ibex/ex_block_i/alu_i/_0841_ ;
 wire \i_ibex/ex_block_i/alu_i/_0842_ ;
 wire \i_ibex/ex_block_i/alu_i/_0843_ ;
 wire \i_ibex/ex_block_i/alu_i/_0844_ ;
 wire net772;
 wire \i_ibex/ex_block_i/alu_i/_0846_ ;
 wire \i_ibex/ex_block_i/alu_i/_0847_ ;
 wire \i_ibex/ex_block_i/alu_i/_0848_ ;
 wire \i_ibex/ex_block_i/alu_i/_0849_ ;
 wire \i_ibex/ex_block_i/alu_i/_0850_ ;
 wire \i_ibex/ex_block_i/alu_i/_0851_ ;
 wire \i_ibex/ex_block_i/alu_i/_0852_ ;
 wire net771;
 wire \i_ibex/ex_block_i/alu_i/_0854_ ;
 wire \i_ibex/ex_block_i/alu_i/_0855_ ;
 wire \i_ibex/ex_block_i/alu_i/_0856_ ;
 wire \i_ibex/ex_block_i/alu_i/_0857_ ;
 wire net770;
 wire \i_ibex/ex_block_i/alu_i/_0859_ ;
 wire \i_ibex/ex_block_i/alu_i/_0860_ ;
 wire \i_ibex/ex_block_i/alu_i/_0861_ ;
 wire \i_ibex/ex_block_i/alu_i/_0862_ ;
 wire \i_ibex/ex_block_i/alu_i/_0863_ ;
 wire \i_ibex/ex_block_i/alu_i/_0864_ ;
 wire \i_ibex/ex_block_i/alu_i/_0865_ ;
 wire \i_ibex/ex_block_i/alu_i/_0866_ ;
 wire \i_ibex/ex_block_i/alu_i/_0867_ ;
 wire \i_ibex/ex_block_i/alu_i/_0868_ ;
 wire net769;
 wire \i_ibex/ex_block_i/alu_i/_0870_ ;
 wire \i_ibex/ex_block_i/alu_i/_0871_ ;
 wire \i_ibex/ex_block_i/alu_i/_0872_ ;
 wire \i_ibex/ex_block_i/alu_i/_0873_ ;
 wire \i_ibex/ex_block_i/alu_i/_0874_ ;
 wire \i_ibex/ex_block_i/alu_i/_0875_ ;
 wire \i_ibex/ex_block_i/alu_i/_0876_ ;
 wire net768;
 wire \i_ibex/ex_block_i/alu_i/_0878_ ;
 wire \i_ibex/ex_block_i/alu_i/_0879_ ;
 wire \i_ibex/ex_block_i/alu_i/_0880_ ;
 wire \i_ibex/ex_block_i/alu_i/_0881_ ;
 wire \i_ibex/ex_block_i/alu_i/_0882_ ;
 wire \i_ibex/ex_block_i/alu_i/_0883_ ;
 wire \i_ibex/ex_block_i/alu_i/_0884_ ;
 wire net767;
 wire \i_ibex/ex_block_i/alu_i/_0886_ ;
 wire \i_ibex/ex_block_i/alu_i/_0887_ ;
 wire \i_ibex/ex_block_i/alu_i/_0888_ ;
 wire \i_ibex/ex_block_i/alu_i/_0889_ ;
 wire net766;
 wire \i_ibex/ex_block_i/alu_i/_0891_ ;
 wire \i_ibex/ex_block_i/alu_i/_0892_ ;
 wire \i_ibex/ex_block_i/alu_i/_0893_ ;
 wire net765;
 wire \i_ibex/ex_block_i/alu_i/_0895_ ;
 wire \i_ibex/ex_block_i/alu_i/_0896_ ;
 wire \i_ibex/ex_block_i/alu_i/_0897_ ;
 wire \i_ibex/ex_block_i/alu_i/_0898_ ;
 wire \i_ibex/ex_block_i/alu_i/_0899_ ;
 wire \i_ibex/ex_block_i/alu_i/_0900_ ;
 wire \i_ibex/ex_block_i/alu_i/_0901_ ;
 wire \i_ibex/ex_block_i/alu_i/_0902_ ;
 wire \i_ibex/ex_block_i/alu_i/_0903_ ;
 wire \i_ibex/ex_block_i/alu_i/_0904_ ;
 wire \i_ibex/ex_block_i/alu_i/_0905_ ;
 wire \i_ibex/ex_block_i/alu_i/_0906_ ;
 wire \i_ibex/ex_block_i/alu_i/_0907_ ;
 wire \i_ibex/ex_block_i/alu_i/_0908_ ;
 wire \i_ibex/ex_block_i/alu_i/_0909_ ;
 wire \i_ibex/ex_block_i/alu_i/_0910_ ;
 wire \i_ibex/ex_block_i/alu_i/_0911_ ;
 wire \i_ibex/ex_block_i/alu_i/_0912_ ;
 wire \i_ibex/ex_block_i/alu_i/_0913_ ;
 wire \i_ibex/ex_block_i/alu_i/_0914_ ;
 wire \i_ibex/ex_block_i/alu_i/_0915_ ;
 wire \i_ibex/ex_block_i/alu_i/_0916_ ;
 wire \i_ibex/ex_block_i/alu_i/_0917_ ;
 wire \i_ibex/ex_block_i/alu_i/_0918_ ;
 wire \i_ibex/ex_block_i/alu_i/_0919_ ;
 wire \i_ibex/ex_block_i/alu_i/_0920_ ;
 wire \i_ibex/ex_block_i/alu_i/_0921_ ;
 wire \i_ibex/ex_block_i/alu_i/_0922_ ;
 wire \i_ibex/ex_block_i/alu_i/_0923_ ;
 wire \i_ibex/ex_block_i/alu_i/_0924_ ;
 wire \i_ibex/ex_block_i/alu_i/_0925_ ;
 wire \i_ibex/ex_block_i/alu_i/_0926_ ;
 wire \i_ibex/ex_block_i/alu_i/_0927_ ;
 wire \i_ibex/ex_block_i/alu_i/_0928_ ;
 wire \i_ibex/ex_block_i/alu_i/_0929_ ;
 wire \i_ibex/ex_block_i/alu_i/_0930_ ;
 wire \i_ibex/ex_block_i/alu_i/_0931_ ;
 wire \i_ibex/ex_block_i/alu_i/_0932_ ;
 wire \i_ibex/ex_block_i/alu_i/_0933_ ;
 wire \i_ibex/ex_block_i/alu_i/_0934_ ;
 wire \i_ibex/ex_block_i/alu_i/_0935_ ;
 wire \i_ibex/ex_block_i/alu_i/_0936_ ;
 wire \i_ibex/ex_block_i/alu_i/_0937_ ;
 wire \i_ibex/ex_block_i/alu_i/_0938_ ;
 wire net764;
 wire \i_ibex/ex_block_i/alu_i/_0940_ ;
 wire \i_ibex/ex_block_i/alu_i/_0941_ ;
 wire \i_ibex/ex_block_i/alu_i/_0942_ ;
 wire \i_ibex/ex_block_i/alu_i/_0943_ ;
 wire \i_ibex/ex_block_i/alu_i/_0944_ ;
 wire \i_ibex/ex_block_i/alu_i/_0945_ ;
 wire \i_ibex/ex_block_i/alu_i/_0946_ ;
 wire \i_ibex/ex_block_i/alu_i/_0947_ ;
 wire \i_ibex/ex_block_i/alu_i/_0948_ ;
 wire \i_ibex/ex_block_i/alu_i/_0949_ ;
 wire \i_ibex/ex_block_i/alu_i/_0950_ ;
 wire \i_ibex/ex_block_i/alu_i/_0951_ ;
 wire \i_ibex/ex_block_i/alu_i/_0952_ ;
 wire \i_ibex/ex_block_i/alu_i/_0953_ ;
 wire \i_ibex/ex_block_i/alu_i/_0954_ ;
 wire \i_ibex/ex_block_i/alu_i/_0955_ ;
 wire \i_ibex/ex_block_i/alu_i/_0956_ ;
 wire \i_ibex/ex_block_i/alu_i/_0957_ ;
 wire \i_ibex/ex_block_i/alu_i/_0958_ ;
 wire \i_ibex/ex_block_i/alu_i/_0959_ ;
 wire \i_ibex/ex_block_i/alu_i/_0960_ ;
 wire \i_ibex/ex_block_i/alu_i/_0961_ ;
 wire \i_ibex/ex_block_i/alu_i/_0962_ ;
 wire \i_ibex/ex_block_i/alu_i/_0963_ ;
 wire \i_ibex/ex_block_i/alu_i/_0964_ ;
 wire \i_ibex/ex_block_i/alu_i/_0965_ ;
 wire \i_ibex/ex_block_i/alu_i/_0966_ ;
 wire \i_ibex/ex_block_i/alu_i/_0967_ ;
 wire \i_ibex/ex_block_i/alu_i/_0968_ ;
 wire \i_ibex/ex_block_i/alu_i/_0969_ ;
 wire \i_ibex/ex_block_i/alu_i/_0970_ ;
 wire \i_ibex/ex_block_i/alu_i/_0971_ ;
 wire \i_ibex/ex_block_i/alu_i/_0972_ ;
 wire net763;
 wire \i_ibex/ex_block_i/alu_i/_0974_ ;
 wire \i_ibex/ex_block_i/alu_i/_0975_ ;
 wire \i_ibex/ex_block_i/alu_i/_0976_ ;
 wire \i_ibex/ex_block_i/alu_i/_0977_ ;
 wire net762;
 wire \i_ibex/ex_block_i/alu_i/_0979_ ;
 wire \i_ibex/ex_block_i/alu_i/_0980_ ;
 wire \i_ibex/ex_block_i/alu_i/_0981_ ;
 wire \i_ibex/ex_block_i/alu_i/_0982_ ;
 wire \i_ibex/ex_block_i/alu_i/_0983_ ;
 wire \i_ibex/ex_block_i/alu_i/_0984_ ;
 wire \i_ibex/ex_block_i/alu_i/_0985_ ;
 wire \i_ibex/ex_block_i/alu_i/_0986_ ;
 wire \i_ibex/ex_block_i/alu_i/_0987_ ;
 wire \i_ibex/ex_block_i/alu_i/_0988_ ;
 wire \i_ibex/ex_block_i/alu_i/_0989_ ;
 wire net761;
 wire \i_ibex/ex_block_i/alu_i/_0991_ ;
 wire \i_ibex/ex_block_i/alu_i/_0992_ ;
 wire \i_ibex/ex_block_i/alu_i/_0993_ ;
 wire \i_ibex/ex_block_i/alu_i/_0994_ ;
 wire \i_ibex/ex_block_i/alu_i/_0995_ ;
 wire \i_ibex/ex_block_i/alu_i/_0996_ ;
 wire \i_ibex/ex_block_i/alu_i/_0997_ ;
 wire net760;
 wire \i_ibex/ex_block_i/alu_i/_0999_ ;
 wire \i_ibex/ex_block_i/alu_i/_1000_ ;
 wire \i_ibex/ex_block_i/alu_i/_1001_ ;
 wire \i_ibex/ex_block_i/alu_i/_1002_ ;
 wire \i_ibex/ex_block_i/alu_i/_1003_ ;
 wire \i_ibex/ex_block_i/alu_i/_1004_ ;
 wire \i_ibex/ex_block_i/alu_i/_1005_ ;
 wire \i_ibex/ex_block_i/alu_i/_1006_ ;
 wire \i_ibex/ex_block_i/alu_i/_1007_ ;
 wire \i_ibex/ex_block_i/alu_i/_1008_ ;
 wire \i_ibex/ex_block_i/alu_i/_1009_ ;
 wire \i_ibex/ex_block_i/alu_i/_1010_ ;
 wire \i_ibex/ex_block_i/alu_i/_1011_ ;
 wire \i_ibex/ex_block_i/alu_i/_1012_ ;
 wire \i_ibex/ex_block_i/alu_i/_1013_ ;
 wire \i_ibex/ex_block_i/alu_i/_1014_ ;
 wire \i_ibex/ex_block_i/alu_i/_1015_ ;
 wire \i_ibex/ex_block_i/alu_i/_1016_ ;
 wire \i_ibex/ex_block_i/alu_i/_1017_ ;
 wire \i_ibex/ex_block_i/alu_i/_1018_ ;
 wire \i_ibex/ex_block_i/alu_i/_1019_ ;
 wire \i_ibex/ex_block_i/alu_i/_1020_ ;
 wire \i_ibex/ex_block_i/alu_i/_1021_ ;
 wire net759;
 wire \i_ibex/ex_block_i/alu_i/_1023_ ;
 wire net758;
 wire \i_ibex/ex_block_i/alu_i/_1025_ ;
 wire \i_ibex/ex_block_i/alu_i/_1026_ ;
 wire \i_ibex/ex_block_i/alu_i/_1027_ ;
 wire \i_ibex/ex_block_i/alu_i/_1028_ ;
 wire \i_ibex/ex_block_i/alu_i/_1029_ ;
 wire \i_ibex/ex_block_i/alu_i/_1030_ ;
 wire \i_ibex/ex_block_i/alu_i/_1031_ ;
 wire \i_ibex/ex_block_i/alu_i/_1032_ ;
 wire \i_ibex/ex_block_i/alu_i/_1033_ ;
 wire \i_ibex/ex_block_i/alu_i/_1034_ ;
 wire \i_ibex/ex_block_i/alu_i/_1035_ ;
 wire \i_ibex/ex_block_i/alu_i/_1036_ ;
 wire \i_ibex/ex_block_i/alu_i/_1037_ ;
 wire \i_ibex/ex_block_i/alu_i/_1038_ ;
 wire net757;
 wire \i_ibex/ex_block_i/alu_i/_1040_ ;
 wire \i_ibex/ex_block_i/alu_i/_1041_ ;
 wire \i_ibex/ex_block_i/alu_i/_1042_ ;
 wire \i_ibex/ex_block_i/alu_i/_1043_ ;
 wire \i_ibex/ex_block_i/alu_i/_1044_ ;
 wire \i_ibex/ex_block_i/alu_i/_1045_ ;
 wire \i_ibex/ex_block_i/alu_i/_1046_ ;
 wire \i_ibex/ex_block_i/alu_i/_1047_ ;
 wire \i_ibex/ex_block_i/alu_i/_1048_ ;
 wire \i_ibex/ex_block_i/alu_i/_1049_ ;
 wire \i_ibex/ex_block_i/alu_i/_1050_ ;
 wire \i_ibex/ex_block_i/alu_i/_1051_ ;
 wire \i_ibex/ex_block_i/alu_i/_1052_ ;
 wire \i_ibex/ex_block_i/alu_i/_1053_ ;
 wire \i_ibex/ex_block_i/alu_i/_1054_ ;
 wire \i_ibex/ex_block_i/alu_i/_1055_ ;
 wire \i_ibex/ex_block_i/alu_i/_1056_ ;
 wire \i_ibex/ex_block_i/alu_i/_1057_ ;
 wire \i_ibex/ex_block_i/alu_i/_1058_ ;
 wire \i_ibex/ex_block_i/alu_i/_1059_ ;
 wire \i_ibex/ex_block_i/alu_i/_1060_ ;
 wire \i_ibex/ex_block_i/alu_i/_1061_ ;
 wire \i_ibex/ex_block_i/alu_i/_1062_ ;
 wire \i_ibex/ex_block_i/alu_i/_1063_ ;
 wire \i_ibex/ex_block_i/alu_i/_1064_ ;
 wire \i_ibex/ex_block_i/alu_i/_1065_ ;
 wire \i_ibex/ex_block_i/alu_i/_1066_ ;
 wire \i_ibex/ex_block_i/alu_i/_1067_ ;
 wire \i_ibex/ex_block_i/alu_i/_1068_ ;
 wire \i_ibex/ex_block_i/alu_i/_1069_ ;
 wire \i_ibex/ex_block_i/alu_i/_1070_ ;
 wire \i_ibex/ex_block_i/alu_i/_1071_ ;
 wire \i_ibex/ex_block_i/alu_i/_1072_ ;
 wire \i_ibex/ex_block_i/alu_i/_1073_ ;
 wire \i_ibex/ex_block_i/alu_i/_1074_ ;
 wire \i_ibex/ex_block_i/alu_i/_1075_ ;
 wire \i_ibex/ex_block_i/alu_i/_1076_ ;
 wire \i_ibex/ex_block_i/alu_i/_1077_ ;
 wire \i_ibex/ex_block_i/alu_i/_1078_ ;
 wire \i_ibex/ex_block_i/alu_i/_1079_ ;
 wire \i_ibex/ex_block_i/alu_i/_1080_ ;
 wire \i_ibex/ex_block_i/alu_i/_1081_ ;
 wire \i_ibex/ex_block_i/alu_i/_1082_ ;
 wire \i_ibex/ex_block_i/alu_i/_1083_ ;
 wire \i_ibex/ex_block_i/alu_i/_1084_ ;
 wire \i_ibex/ex_block_i/alu_i/_1085_ ;
 wire \i_ibex/ex_block_i/alu_i/_1086_ ;
 wire \i_ibex/ex_block_i/alu_i/_1087_ ;
 wire \i_ibex/ex_block_i/alu_i/_1088_ ;
 wire \i_ibex/ex_block_i/alu_i/_1089_ ;
 wire \i_ibex/ex_block_i/alu_i/_1090_ ;
 wire \i_ibex/ex_block_i/alu_i/_1091_ ;
 wire \i_ibex/ex_block_i/alu_i/_1092_ ;
 wire net756;
 wire net755;
 wire net754;
 wire net753;
 wire \i_ibex/ex_block_i/alu_i/_1097_ ;
 wire \i_ibex/ex_block_i/alu_i/_1098_ ;
 wire \i_ibex/ex_block_i/alu_i/_1099_ ;
 wire net752;
 wire \i_ibex/ex_block_i/alu_i/_1101_ ;
 wire \i_ibex/ex_block_i/alu_i/_1102_ ;
 wire \i_ibex/ex_block_i/alu_i/_1103_ ;
 wire \i_ibex/ex_block_i/alu_i/_1104_ ;
 wire \i_ibex/ex_block_i/alu_i/_1105_ ;
 wire \i_ibex/ex_block_i/alu_i/_1106_ ;
 wire \i_ibex/ex_block_i/alu_i/_1107_ ;
 wire \i_ibex/ex_block_i/alu_i/_1108_ ;
 wire \i_ibex/ex_block_i/alu_i/_1109_ ;
 wire \i_ibex/ex_block_i/alu_i/_1110_ ;
 wire \i_ibex/ex_block_i/alu_i/_1111_ ;
 wire net751;
 wire \i_ibex/ex_block_i/alu_i/_1113_ ;
 wire \i_ibex/ex_block_i/alu_i/_1114_ ;
 wire \i_ibex/ex_block_i/alu_i/_1115_ ;
 wire \i_ibex/ex_block_i/alu_i/_1116_ ;
 wire \i_ibex/ex_block_i/alu_i/_1117_ ;
 wire \i_ibex/ex_block_i/alu_i/_1118_ ;
 wire \i_ibex/ex_block_i/alu_i/_1119_ ;
 wire net750;
 wire \i_ibex/ex_block_i/alu_i/_1121_ ;
 wire \i_ibex/ex_block_i/alu_i/_1122_ ;
 wire \i_ibex/ex_block_i/alu_i/_1123_ ;
 wire \i_ibex/ex_block_i/alu_i/_1124_ ;
 wire \i_ibex/ex_block_i/alu_i/_1125_ ;
 wire \i_ibex/ex_block_i/alu_i/_1126_ ;
 wire \i_ibex/ex_block_i/alu_i/_1127_ ;
 wire \i_ibex/ex_block_i/alu_i/_1128_ ;
 wire \i_ibex/ex_block_i/alu_i/_1129_ ;
 wire \i_ibex/ex_block_i/alu_i/_1130_ ;
 wire \i_ibex/ex_block_i/alu_i/_1131_ ;
 wire \i_ibex/ex_block_i/alu_i/_1132_ ;
 wire \i_ibex/ex_block_i/alu_i/_1133_ ;
 wire \i_ibex/ex_block_i/alu_i/_1134_ ;
 wire \i_ibex/ex_block_i/alu_i/_1135_ ;
 wire \i_ibex/ex_block_i/alu_i/_1136_ ;
 wire \i_ibex/ex_block_i/alu_i/_1137_ ;
 wire \i_ibex/ex_block_i/alu_i/_1138_ ;
 wire \i_ibex/ex_block_i/alu_i/_1139_ ;
 wire \i_ibex/ex_block_i/alu_i/_1140_ ;
 wire net749;
 wire \i_ibex/ex_block_i/alu_i/_1142_ ;
 wire \i_ibex/ex_block_i/alu_i/_1143_ ;
 wire \i_ibex/ex_block_i/alu_i/_1144_ ;
 wire \i_ibex/ex_block_i/alu_i/_1145_ ;
 wire \i_ibex/ex_block_i/alu_i/_1146_ ;
 wire \i_ibex/ex_block_i/alu_i/_1147_ ;
 wire \i_ibex/ex_block_i/alu_i/_1148_ ;
 wire \i_ibex/ex_block_i/alu_i/_1149_ ;
 wire \i_ibex/ex_block_i/alu_i/_1150_ ;
 wire net748;
 wire \i_ibex/ex_block_i/alu_i/_1152_ ;
 wire \i_ibex/ex_block_i/alu_i/_1153_ ;
 wire \i_ibex/ex_block_i/alu_i/_1154_ ;
 wire \i_ibex/ex_block_i/alu_i/_1155_ ;
 wire \i_ibex/ex_block_i/alu_i/_1156_ ;
 wire \i_ibex/ex_block_i/alu_i/_1157_ ;
 wire \i_ibex/ex_block_i/alu_i/_1158_ ;
 wire \i_ibex/ex_block_i/alu_i/_1159_ ;
 wire \i_ibex/ex_block_i/alu_i/_1160_ ;
 wire \i_ibex/ex_block_i/alu_i/_1161_ ;
 wire \i_ibex/ex_block_i/alu_i/_1162_ ;
 wire \i_ibex/ex_block_i/alu_i/_1163_ ;
 wire \i_ibex/ex_block_i/alu_i/_1164_ ;
 wire \i_ibex/ex_block_i/alu_i/_1165_ ;
 wire \i_ibex/ex_block_i/alu_i/_1166_ ;
 wire \i_ibex/ex_block_i/alu_i/_1167_ ;
 wire \i_ibex/ex_block_i/alu_i/_1168_ ;
 wire \i_ibex/ex_block_i/alu_i/_1169_ ;
 wire \i_ibex/ex_block_i/alu_i/_1170_ ;
 wire \i_ibex/ex_block_i/alu_i/_1171_ ;
 wire \i_ibex/ex_block_i/alu_i/_1172_ ;
 wire \i_ibex/ex_block_i/alu_i/_1173_ ;
 wire \i_ibex/ex_block_i/alu_i/_1174_ ;
 wire \i_ibex/ex_block_i/alu_i/_1175_ ;
 wire \i_ibex/ex_block_i/alu_i/_1176_ ;
 wire \i_ibex/ex_block_i/alu_i/_1177_ ;
 wire \i_ibex/ex_block_i/alu_i/_1178_ ;
 wire \i_ibex/ex_block_i/alu_i/_1179_ ;
 wire \i_ibex/ex_block_i/alu_i/_1180_ ;
 wire \i_ibex/ex_block_i/alu_i/_1181_ ;
 wire \i_ibex/ex_block_i/alu_i/_1182_ ;
 wire \i_ibex/ex_block_i/alu_i/_1183_ ;
 wire \i_ibex/ex_block_i/alu_i/_1184_ ;
 wire \i_ibex/ex_block_i/alu_i/_1185_ ;
 wire \i_ibex/ex_block_i/alu_i/_1186_ ;
 wire \i_ibex/ex_block_i/alu_i/_1187_ ;
 wire \i_ibex/ex_block_i/alu_i/_1188_ ;
 wire \i_ibex/ex_block_i/alu_i/_1189_ ;
 wire \i_ibex/ex_block_i/alu_i/_1190_ ;
 wire \i_ibex/ex_block_i/alu_i/_1191_ ;
 wire \i_ibex/ex_block_i/alu_i/_1192_ ;
 wire \i_ibex/ex_block_i/alu_i/_1193_ ;
 wire \i_ibex/ex_block_i/alu_i/_1194_ ;
 wire \i_ibex/ex_block_i/alu_i/_1195_ ;
 wire \i_ibex/ex_block_i/alu_i/_1196_ ;
 wire \i_ibex/ex_block_i/alu_i/_1197_ ;
 wire \i_ibex/ex_block_i/alu_i/_1198_ ;
 wire \i_ibex/ex_block_i/alu_i/_1199_ ;
 wire \i_ibex/ex_block_i/alu_i/_1200_ ;
 wire \i_ibex/ex_block_i/alu_i/_1201_ ;
 wire \i_ibex/ex_block_i/alu_i/_1202_ ;
 wire \i_ibex/ex_block_i/alu_i/_1203_ ;
 wire \i_ibex/ex_block_i/alu_i/_1204_ ;
 wire \i_ibex/ex_block_i/alu_i/_1205_ ;
 wire \i_ibex/ex_block_i/alu_i/_1206_ ;
 wire \i_ibex/ex_block_i/alu_i/_1207_ ;
 wire \i_ibex/ex_block_i/alu_i/_1208_ ;
 wire \i_ibex/ex_block_i/alu_i/_1209_ ;
 wire \i_ibex/ex_block_i/alu_i/_1210_ ;
 wire \i_ibex/ex_block_i/alu_i/_1211_ ;
 wire \i_ibex/ex_block_i/alu_i/_1212_ ;
 wire \i_ibex/ex_block_i/alu_i/_1213_ ;
 wire \i_ibex/ex_block_i/alu_i/_1214_ ;
 wire \i_ibex/ex_block_i/alu_i/_1215_ ;
 wire \i_ibex/ex_block_i/alu_i/_1216_ ;
 wire \i_ibex/ex_block_i/alu_i/_1217_ ;
 wire \i_ibex/ex_block_i/alu_i/_1218_ ;
 wire \i_ibex/ex_block_i/alu_i/_1219_ ;
 wire \i_ibex/ex_block_i/alu_i/_1220_ ;
 wire \i_ibex/ex_block_i/alu_i/_1221_ ;
 wire \i_ibex/ex_block_i/alu_i/_1222_ ;
 wire \i_ibex/ex_block_i/alu_i/_1223_ ;
 wire \i_ibex/ex_block_i/alu_i/_1224_ ;
 wire \i_ibex/ex_block_i/alu_i/_1225_ ;
 wire \i_ibex/ex_block_i/alu_i/_1226_ ;
 wire \i_ibex/ex_block_i/alu_i/_1227_ ;
 wire \i_ibex/ex_block_i/alu_i/_1228_ ;
 wire \i_ibex/ex_block_i/alu_i/_1229_ ;
 wire \i_ibex/ex_block_i/alu_i/_1230_ ;
 wire \i_ibex/ex_block_i/alu_i/_1231_ ;
 wire \i_ibex/ex_block_i/alu_i/_1232_ ;
 wire \i_ibex/ex_block_i/alu_i/_1233_ ;
 wire \i_ibex/ex_block_i/alu_i/_1234_ ;
 wire \i_ibex/ex_block_i/alu_i/_1235_ ;
 wire \i_ibex/ex_block_i/alu_i/_1236_ ;
 wire \i_ibex/ex_block_i/alu_i/_1237_ ;
 wire \i_ibex/ex_block_i/alu_i/_1238_ ;
 wire \i_ibex/ex_block_i/alu_i/_1239_ ;
 wire \i_ibex/ex_block_i/alu_i/_1240_ ;
 wire \i_ibex/ex_block_i/alu_i/_1241_ ;
 wire \i_ibex/ex_block_i/alu_i/_1242_ ;
 wire \i_ibex/ex_block_i/alu_i/_1243_ ;
 wire \i_ibex/ex_block_i/alu_i/_1244_ ;
 wire \i_ibex/ex_block_i/alu_i/_1245_ ;
 wire \i_ibex/ex_block_i/alu_i/_1246_ ;
 wire \i_ibex/ex_block_i/alu_i/_1247_ ;
 wire \i_ibex/ex_block_i/alu_i/_1248_ ;
 wire \i_ibex/ex_block_i/alu_i/_1249_ ;
 wire \i_ibex/ex_block_i/alu_i/_1250_ ;
 wire \i_ibex/ex_block_i/alu_i/_1251_ ;
 wire \i_ibex/ex_block_i/alu_i/_1252_ ;
 wire \i_ibex/ex_block_i/alu_i/_1253_ ;
 wire \i_ibex/ex_block_i/alu_i/_1254_ ;
 wire \i_ibex/ex_block_i/alu_i/_1255_ ;
 wire \i_ibex/ex_block_i/alu_i/_1256_ ;
 wire \i_ibex/ex_block_i/alu_i/_1257_ ;
 wire \i_ibex/ex_block_i/alu_i/_1258_ ;
 wire \i_ibex/ex_block_i/alu_i/_1259_ ;
 wire \i_ibex/ex_block_i/alu_i/_1260_ ;
 wire \i_ibex/ex_block_i/alu_i/_1261_ ;
 wire \i_ibex/ex_block_i/alu_i/_1262_ ;
 wire \i_ibex/ex_block_i/alu_i/_1263_ ;
 wire \i_ibex/ex_block_i/alu_i/_1264_ ;
 wire net747;
 wire \i_ibex/ex_block_i/alu_i/_1266_ ;
 wire \i_ibex/ex_block_i/alu_i/_1267_ ;
 wire \i_ibex/ex_block_i/alu_i/_1268_ ;
 wire \i_ibex/ex_block_i/alu_i/_1269_ ;
 wire \i_ibex/ex_block_i/alu_i/_1270_ ;
 wire \i_ibex/ex_block_i/alu_i/_1271_ ;
 wire \i_ibex/ex_block_i/alu_i/_1272_ ;
 wire \i_ibex/ex_block_i/alu_i/_1273_ ;
 wire net746;
 wire \i_ibex/ex_block_i/alu_i/_1275_ ;
 wire \i_ibex/ex_block_i/alu_i/_1276_ ;
 wire \i_ibex/ex_block_i/alu_i/_1277_ ;
 wire \i_ibex/ex_block_i/alu_i/_1278_ ;
 wire \i_ibex/ex_block_i/alu_i/_1279_ ;
 wire \i_ibex/ex_block_i/alu_i/_1280_ ;
 wire \i_ibex/ex_block_i/alu_i/_1281_ ;
 wire \i_ibex/ex_block_i/alu_i/_1282_ ;
 wire \i_ibex/ex_block_i/alu_i/_1283_ ;
 wire \i_ibex/ex_block_i/alu_i/_1284_ ;
 wire \i_ibex/ex_block_i/alu_i/_1285_ ;
 wire \i_ibex/ex_block_i/alu_i/_1286_ ;
 wire \i_ibex/ex_block_i/alu_i/_1287_ ;
 wire net745;
 wire \i_ibex/ex_block_i/alu_i/_1289_ ;
 wire \i_ibex/ex_block_i/alu_i/_1290_ ;
 wire \i_ibex/ex_block_i/alu_i/_1291_ ;
 wire \i_ibex/ex_block_i/alu_i/_1292_ ;
 wire \i_ibex/ex_block_i/alu_i/_1293_ ;
 wire \i_ibex/ex_block_i/alu_i/_1294_ ;
 wire \i_ibex/ex_block_i/alu_i/_1295_ ;
 wire \i_ibex/ex_block_i/alu_i/_1296_ ;
 wire \i_ibex/ex_block_i/alu_i/_1297_ ;
 wire \i_ibex/ex_block_i/alu_i/_1298_ ;
 wire \i_ibex/ex_block_i/alu_i/_1299_ ;
 wire \i_ibex/ex_block_i/alu_i/_1300_ ;
 wire \i_ibex/ex_block_i/alu_i/_1301_ ;
 wire \i_ibex/ex_block_i/alu_i/_1302_ ;
 wire \i_ibex/ex_block_i/alu_i/_1303_ ;
 wire \i_ibex/ex_block_i/alu_i/_1304_ ;
 wire \i_ibex/ex_block_i/alu_i/_1305_ ;
 wire \i_ibex/ex_block_i/alu_i/_1306_ ;
 wire \i_ibex/ex_block_i/alu_i/_1307_ ;
 wire \i_ibex/ex_block_i/alu_i/_1308_ ;
 wire \i_ibex/ex_block_i/alu_i/_1309_ ;
 wire \i_ibex/ex_block_i/alu_i/_1310_ ;
 wire \i_ibex/ex_block_i/alu_i/_1311_ ;
 wire \i_ibex/ex_block_i/alu_i/_1312_ ;
 wire \i_ibex/ex_block_i/alu_i/_1313_ ;
 wire \i_ibex/ex_block_i/alu_i/_1314_ ;
 wire \i_ibex/ex_block_i/alu_i/_1315_ ;
 wire \i_ibex/ex_block_i/alu_i/_1316_ ;
 wire \i_ibex/ex_block_i/alu_i/_1317_ ;
 wire \i_ibex/ex_block_i/alu_i/_1318_ ;
 wire \i_ibex/ex_block_i/alu_i/_1319_ ;
 wire \i_ibex/ex_block_i/alu_i/_1320_ ;
 wire \i_ibex/ex_block_i/alu_i/_1321_ ;
 wire \i_ibex/ex_block_i/alu_i/_1322_ ;
 wire \i_ibex/ex_block_i/alu_i/_1323_ ;
 wire \i_ibex/ex_block_i/alu_i/_1324_ ;
 wire \i_ibex/ex_block_i/alu_i/_1325_ ;
 wire \i_ibex/ex_block_i/alu_i/_1326_ ;
 wire \i_ibex/ex_block_i/alu_i/_1327_ ;
 wire \i_ibex/ex_block_i/alu_i/_1328_ ;
 wire \i_ibex/ex_block_i/alu_i/_1329_ ;
 wire \i_ibex/ex_block_i/alu_i/_1330_ ;
 wire \i_ibex/ex_block_i/alu_i/_1331_ ;
 wire \i_ibex/ex_block_i/alu_i/_1332_ ;
 wire \i_ibex/ex_block_i/alu_i/_1333_ ;
 wire \i_ibex/ex_block_i/alu_i/_1334_ ;
 wire \i_ibex/ex_block_i/alu_i/_1335_ ;
 wire \i_ibex/ex_block_i/alu_i/_1336_ ;
 wire \i_ibex/ex_block_i/alu_i/_1337_ ;
 wire \i_ibex/ex_block_i/alu_i/_1338_ ;
 wire \i_ibex/ex_block_i/alu_i/_1339_ ;
 wire \i_ibex/ex_block_i/alu_i/_1340_ ;
 wire \i_ibex/ex_block_i/alu_i/_1341_ ;
 wire \i_ibex/ex_block_i/alu_i/_1342_ ;
 wire \i_ibex/ex_block_i/alu_i/_1343_ ;
 wire \i_ibex/ex_block_i/alu_i/_1344_ ;
 wire \i_ibex/ex_block_i/alu_i/_1345_ ;
 wire \i_ibex/ex_block_i/alu_i/_1346_ ;
 wire \i_ibex/ex_block_i/alu_i/_1347_ ;
 wire \i_ibex/id_stage_i/_0000_ ;
 wire \i_ibex/id_stage_i/_0001_ ;
 wire \i_ibex/id_stage_i/_0002_ ;
 wire \i_ibex/id_stage_i/_0003_ ;
 wire \i_ibex/id_stage_i/_0004_ ;
 wire \i_ibex/id_stage_i/_0005_ ;
 wire \i_ibex/id_stage_i/_0006_ ;
 wire \i_ibex/id_stage_i/_0007_ ;
 wire \i_ibex/id_stage_i/_0008_ ;
 wire \i_ibex/id_stage_i/_0009_ ;
 wire \i_ibex/id_stage_i/_0010_ ;
 wire \i_ibex/id_stage_i/_0011_ ;
 wire \i_ibex/id_stage_i/_0012_ ;
 wire \i_ibex/id_stage_i/_0013_ ;
 wire \i_ibex/id_stage_i/_0014_ ;
 wire \i_ibex/id_stage_i/_0015_ ;
 wire \i_ibex/id_stage_i/_0016_ ;
 wire \i_ibex/id_stage_i/_0017_ ;
 wire \i_ibex/id_stage_i/_0018_ ;
 wire \i_ibex/id_stage_i/_0019_ ;
 wire \i_ibex/id_stage_i/_0020_ ;
 wire \i_ibex/id_stage_i/_0021_ ;
 wire \i_ibex/id_stage_i/_0022_ ;
 wire \i_ibex/id_stage_i/_0023_ ;
 wire \i_ibex/id_stage_i/_0024_ ;
 wire \i_ibex/id_stage_i/_0025_ ;
 wire \i_ibex/id_stage_i/_0026_ ;
 wire \i_ibex/id_stage_i/_0027_ ;
 wire \i_ibex/id_stage_i/_0028_ ;
 wire \i_ibex/id_stage_i/_0029_ ;
 wire \i_ibex/id_stage_i/_0030_ ;
 wire \i_ibex/id_stage_i/_0031_ ;
 wire \i_ibex/id_stage_i/_0032_ ;
 wire \i_ibex/id_stage_i/_0033_ ;
 wire \i_ibex/id_stage_i/_0034_ ;
 wire \i_ibex/id_stage_i/_0035_ ;
 wire \i_ibex/id_stage_i/_0036_ ;
 wire \i_ibex/id_stage_i/_0037_ ;
 wire \i_ibex/id_stage_i/_0038_ ;
 wire \i_ibex/id_stage_i/_0039_ ;
 wire \i_ibex/id_stage_i/_0040_ ;
 wire \i_ibex/id_stage_i/_0041_ ;
 wire \i_ibex/id_stage_i/_0042_ ;
 wire \i_ibex/id_stage_i/_0043_ ;
 wire \i_ibex/id_stage_i/_0044_ ;
 wire \i_ibex/id_stage_i/_0045_ ;
 wire \i_ibex/id_stage_i/_0046_ ;
 wire \i_ibex/id_stage_i/_0047_ ;
 wire \i_ibex/id_stage_i/_0048_ ;
 wire \i_ibex/id_stage_i/_0049_ ;
 wire \i_ibex/id_stage_i/_0050_ ;
 wire \i_ibex/id_stage_i/_0051_ ;
 wire \i_ibex/id_stage_i/_0052_ ;
 wire \i_ibex/id_stage_i/_0053_ ;
 wire \i_ibex/id_stage_i/_0054_ ;
 wire \i_ibex/id_stage_i/_0055_ ;
 wire \i_ibex/id_stage_i/_0056_ ;
 wire \i_ibex/id_stage_i/_0057_ ;
 wire \i_ibex/id_stage_i/_0058_ ;
 wire \i_ibex/id_stage_i/_0059_ ;
 wire \i_ibex/id_stage_i/_0060_ ;
 wire \i_ibex/id_stage_i/_0061_ ;
 wire \i_ibex/id_stage_i/_0062_ ;
 wire \i_ibex/id_stage_i/_0063_ ;
 wire \i_ibex/id_stage_i/_0064_ ;
 wire \i_ibex/id_stage_i/_0065_ ;
 wire \i_ibex/id_stage_i/_0066_ ;
 wire \i_ibex/id_stage_i/_0067_ ;
 wire \i_ibex/id_stage_i/_0068_ ;
 wire \i_ibex/id_stage_i/_0069_ ;
 wire \i_ibex/id_stage_i/_0070_ ;
 wire \i_ibex/id_stage_i/_0071_ ;
 wire \i_ibex/id_stage_i/_0072_ ;
 wire \i_ibex/id_stage_i/_0073_ ;
 wire \i_ibex/id_stage_i/_0074_ ;
 wire \i_ibex/id_stage_i/_0075_ ;
 wire \i_ibex/id_stage_i/_0076_ ;
 wire \i_ibex/id_stage_i/_0077_ ;
 wire \i_ibex/id_stage_i/_0078_ ;
 wire \i_ibex/id_stage_i/_0079_ ;
 wire \i_ibex/id_stage_i/_0080_ ;
 wire \i_ibex/id_stage_i/_0081_ ;
 wire net651;
 wire \i_ibex/id_stage_i/_0083_ ;
 wire \i_ibex/id_stage_i/_0084_ ;
 wire \i_ibex/id_stage_i/_0085_ ;
 wire \i_ibex/id_stage_i/_0086_ ;
 wire \i_ibex/id_stage_i/_0087_ ;
 wire \i_ibex/id_stage_i/_0088_ ;
 wire \i_ibex/id_stage_i/_0089_ ;
 wire \i_ibex/id_stage_i/_0090_ ;
 wire \i_ibex/id_stage_i/_0091_ ;
 wire \i_ibex/id_stage_i/_0092_ ;
 wire \i_ibex/id_stage_i/_0093_ ;
 wire \i_ibex/id_stage_i/_0094_ ;
 wire \i_ibex/id_stage_i/_0095_ ;
 wire net650;
 wire \i_ibex/id_stage_i/_0097_ ;
 wire \i_ibex/id_stage_i/_0098_ ;
 wire \i_ibex/id_stage_i/_0099_ ;
 wire \i_ibex/id_stage_i/_0100_ ;
 wire \i_ibex/id_stage_i/_0101_ ;
 wire \i_ibex/id_stage_i/_0102_ ;
 wire net649;
 wire \i_ibex/id_stage_i/_0104_ ;
 wire \i_ibex/id_stage_i/_0105_ ;
 wire \i_ibex/id_stage_i/_0106_ ;
 wire \i_ibex/id_stage_i/_0107_ ;
 wire \i_ibex/id_stage_i/_0108_ ;
 wire \i_ibex/id_stage_i/_0109_ ;
 wire net648;
 wire \i_ibex/id_stage_i/_0111_ ;
 wire \i_ibex/id_stage_i/_0112_ ;
 wire \i_ibex/id_stage_i/_0113_ ;
 wire \i_ibex/id_stage_i/_0114_ ;
 wire \i_ibex/id_stage_i/_0115_ ;
 wire \i_ibex/id_stage_i/_0116_ ;
 wire \i_ibex/id_stage_i/_0117_ ;
 wire net647;
 wire \i_ibex/id_stage_i/_0119_ ;
 wire \i_ibex/id_stage_i/_0120_ ;
 wire net646;
 wire \i_ibex/id_stage_i/_0122_ ;
 wire \i_ibex/id_stage_i/_0123_ ;
 wire \i_ibex/id_stage_i/_0124_ ;
 wire net645;
 wire \i_ibex/id_stage_i/_0126_ ;
 wire \i_ibex/id_stage_i/_0127_ ;
 wire \i_ibex/id_stage_i/_0128_ ;
 wire net644;
 wire \i_ibex/id_stage_i/_0130_ ;
 wire \i_ibex/id_stage_i/_0131_ ;
 wire net643;
 wire \i_ibex/id_stage_i/_0133_ ;
 wire \i_ibex/id_stage_i/_0134_ ;
 wire \i_ibex/id_stage_i/_0135_ ;
 wire \i_ibex/id_stage_i/_0136_ ;
 wire \i_ibex/id_stage_i/_0137_ ;
 wire \i_ibex/id_stage_i/_0138_ ;
 wire \i_ibex/id_stage_i/_0139_ ;
 wire net642;
 wire \i_ibex/id_stage_i/_0141_ ;
 wire \i_ibex/id_stage_i/_0142_ ;
 wire \i_ibex/id_stage_i/_0143_ ;
 wire \i_ibex/id_stage_i/_0144_ ;
 wire \i_ibex/id_stage_i/_0145_ ;
 wire \i_ibex/id_stage_i/_0146_ ;
 wire \i_ibex/id_stage_i/_0147_ ;
 wire \i_ibex/id_stage_i/_0148_ ;
 wire \i_ibex/id_stage_i/_0149_ ;
 wire \i_ibex/id_stage_i/_0150_ ;
 wire \i_ibex/id_stage_i/_0151_ ;
 wire \i_ibex/id_stage_i/_0152_ ;
 wire \i_ibex/id_stage_i/_0153_ ;
 wire \i_ibex/id_stage_i/_0154_ ;
 wire \i_ibex/id_stage_i/_0155_ ;
 wire \i_ibex/id_stage_i/_0156_ ;
 wire \i_ibex/id_stage_i/_0157_ ;
 wire \i_ibex/id_stage_i/_0158_ ;
 wire \i_ibex/id_stage_i/_0159_ ;
 wire \i_ibex/id_stage_i/_0160_ ;
 wire \i_ibex/id_stage_i/_0161_ ;
 wire \i_ibex/id_stage_i/_0162_ ;
 wire net641;
 wire \i_ibex/id_stage_i/_0164_ ;
 wire \i_ibex/id_stage_i/_0165_ ;
 wire \i_ibex/id_stage_i/_0166_ ;
 wire \i_ibex/id_stage_i/_0167_ ;
 wire \i_ibex/id_stage_i/_0168_ ;
 wire \i_ibex/id_stage_i/_0169_ ;
 wire \i_ibex/id_stage_i/_0170_ ;
 wire \i_ibex/id_stage_i/_0171_ ;
 wire \i_ibex/id_stage_i/_0172_ ;
 wire \i_ibex/id_stage_i/_0173_ ;
 wire \i_ibex/id_stage_i/_0174_ ;
 wire \i_ibex/id_stage_i/_0175_ ;
 wire net640;
 wire \i_ibex/id_stage_i/_0177_ ;
 wire \i_ibex/id_stage_i/_0178_ ;
 wire \i_ibex/id_stage_i/_0179_ ;
 wire \i_ibex/id_stage_i/_0180_ ;
 wire \i_ibex/id_stage_i/_0181_ ;
 wire \i_ibex/id_stage_i/_0182_ ;
 wire net639;
 wire \i_ibex/id_stage_i/_0184_ ;
 wire \i_ibex/id_stage_i/_0185_ ;
 wire \i_ibex/id_stage_i/_0186_ ;
 wire \i_ibex/id_stage_i/_0187_ ;
 wire \i_ibex/id_stage_i/_0188_ ;
 wire \i_ibex/id_stage_i/_0189_ ;
 wire net638;
 wire \i_ibex/id_stage_i/_0191_ ;
 wire \i_ibex/id_stage_i/_0192_ ;
 wire \i_ibex/id_stage_i/_0193_ ;
 wire \i_ibex/id_stage_i/_0194_ ;
 wire \i_ibex/id_stage_i/_0195_ ;
 wire \i_ibex/id_stage_i/_0196_ ;
 wire \i_ibex/id_stage_i/_0197_ ;
 wire net637;
 wire \i_ibex/id_stage_i/_0199_ ;
 wire \i_ibex/id_stage_i/_0200_ ;
 wire net636;
 wire \i_ibex/id_stage_i/_0202_ ;
 wire \i_ibex/id_stage_i/_0203_ ;
 wire \i_ibex/id_stage_i/_0204_ ;
 wire net635;
 wire \i_ibex/id_stage_i/_0206_ ;
 wire \i_ibex/id_stage_i/_0207_ ;
 wire \i_ibex/id_stage_i/_0208_ ;
 wire net634;
 wire \i_ibex/id_stage_i/_0210_ ;
 wire \i_ibex/id_stage_i/_0211_ ;
 wire \i_ibex/id_stage_i/_0212_ ;
 wire \i_ibex/id_stage_i/_0213_ ;
 wire \i_ibex/id_stage_i/_0214_ ;
 wire \i_ibex/id_stage_i/_0215_ ;
 wire \i_ibex/id_stage_i/_0216_ ;
 wire \i_ibex/id_stage_i/_0217_ ;
 wire \i_ibex/id_stage_i/_0218_ ;
 wire \i_ibex/id_stage_i/_0219_ ;
 wire \i_ibex/id_stage_i/_0220_ ;
 wire \i_ibex/id_stage_i/_0221_ ;
 wire \i_ibex/id_stage_i/_0222_ ;
 wire \i_ibex/id_stage_i/_0223_ ;
 wire \i_ibex/id_stage_i/_0224_ ;
 wire \i_ibex/id_stage_i/_0225_ ;
 wire \i_ibex/id_stage_i/_0226_ ;
 wire \i_ibex/id_stage_i/_0227_ ;
 wire \i_ibex/id_stage_i/_0228_ ;
 wire \i_ibex/id_stage_i/_0229_ ;
 wire \i_ibex/id_stage_i/_0230_ ;
 wire \i_ibex/id_stage_i/_0231_ ;
 wire \i_ibex/id_stage_i/_0232_ ;
 wire \i_ibex/id_stage_i/_0233_ ;
 wire \i_ibex/id_stage_i/_0234_ ;
 wire \i_ibex/id_stage_i/_0235_ ;
 wire \i_ibex/id_stage_i/_0236_ ;
 wire \i_ibex/id_stage_i/_0237_ ;
 wire \i_ibex/id_stage_i/_0238_ ;
 wire \i_ibex/id_stage_i/_0239_ ;
 wire \i_ibex/id_stage_i/_0240_ ;
 wire \i_ibex/id_stage_i/_0241_ ;
 wire \i_ibex/id_stage_i/_0242_ ;
 wire \i_ibex/id_stage_i/_0243_ ;
 wire \i_ibex/id_stage_i/_0244_ ;
 wire \i_ibex/id_stage_i/_0245_ ;
 wire \i_ibex/id_stage_i/_0246_ ;
 wire \i_ibex/id_stage_i/_0247_ ;
 wire \i_ibex/id_stage_i/_0248_ ;
 wire \i_ibex/id_stage_i/_0249_ ;
 wire \i_ibex/id_stage_i/_0250_ ;
 wire \i_ibex/id_stage_i/_0251_ ;
 wire \i_ibex/id_stage_i/_0252_ ;
 wire \i_ibex/id_stage_i/_0253_ ;
 wire \i_ibex/id_stage_i/_0254_ ;
 wire \i_ibex/id_stage_i/_0255_ ;
 wire \i_ibex/id_stage_i/_0256_ ;
 wire \i_ibex/id_stage_i/_0257_ ;
 wire \i_ibex/id_stage_i/_0258_ ;
 wire \i_ibex/id_stage_i/_0259_ ;
 wire \i_ibex/id_stage_i/_0260_ ;
 wire \i_ibex/id_stage_i/_0261_ ;
 wire \i_ibex/id_stage_i/_0262_ ;
 wire \i_ibex/id_stage_i/_0263_ ;
 wire \i_ibex/id_stage_i/_0264_ ;
 wire \i_ibex/id_stage_i/_0265_ ;
 wire \i_ibex/id_stage_i/_0266_ ;
 wire \i_ibex/id_stage_i/_0267_ ;
 wire \i_ibex/id_stage_i/_0268_ ;
 wire \i_ibex/id_stage_i/_0269_ ;
 wire \i_ibex/id_stage_i/_0270_ ;
 wire \i_ibex/id_stage_i/_0271_ ;
 wire \i_ibex/id_stage_i/_0272_ ;
 wire \i_ibex/id_stage_i/_0273_ ;
 wire \i_ibex/id_stage_i/_0274_ ;
 wire \i_ibex/id_stage_i/_0275_ ;
 wire \i_ibex/id_stage_i/_0276_ ;
 wire \i_ibex/id_stage_i/_0277_ ;
 wire \i_ibex/id_stage_i/_0278_ ;
 wire \i_ibex/id_stage_i/_0279_ ;
 wire \i_ibex/id_stage_i/_0280_ ;
 wire \i_ibex/id_stage_i/_0281_ ;
 wire \i_ibex/id_stage_i/_0282_ ;
 wire \i_ibex/id_stage_i/_0283_ ;
 wire \i_ibex/id_stage_i/_0284_ ;
 wire \i_ibex/id_stage_i/_0285_ ;
 wire \i_ibex/id_stage_i/_0286_ ;
 wire \i_ibex/id_stage_i/_0287_ ;
 wire \i_ibex/id_stage_i/_0288_ ;
 wire \i_ibex/id_stage_i/_0289_ ;
 wire \i_ibex/id_stage_i/_0290_ ;
 wire \i_ibex/id_stage_i/_0291_ ;
 wire \i_ibex/id_stage_i/_0292_ ;
 wire \i_ibex/id_stage_i/_0293_ ;
 wire \i_ibex/id_stage_i/_0294_ ;
 wire \i_ibex/id_stage_i/_0295_ ;
 wire \i_ibex/id_stage_i/_0296_ ;
 wire \i_ibex/id_stage_i/_0297_ ;
 wire \i_ibex/id_stage_i/_0298_ ;
 wire \i_ibex/id_stage_i/_0299_ ;
 wire \i_ibex/id_stage_i/_0300_ ;
 wire \i_ibex/id_stage_i/_0301_ ;
 wire \i_ibex/id_stage_i/_0302_ ;
 wire \i_ibex/id_stage_i/_0303_ ;
 wire \i_ibex/id_stage_i/_0304_ ;
 wire \i_ibex/id_stage_i/_0305_ ;
 wire \i_ibex/id_stage_i/_0306_ ;
 wire \i_ibex/id_stage_i/_0307_ ;
 wire \i_ibex/id_stage_i/_0308_ ;
 wire \i_ibex/id_stage_i/_0309_ ;
 wire \i_ibex/id_stage_i/_0310_ ;
 wire \i_ibex/id_stage_i/_0311_ ;
 wire \i_ibex/id_stage_i/_0312_ ;
 wire \i_ibex/id_stage_i/_0313_ ;
 wire \i_ibex/id_stage_i/_0314_ ;
 wire \i_ibex/id_stage_i/_0315_ ;
 wire \i_ibex/id_stage_i/_0316_ ;
 wire \i_ibex/id_stage_i/_0317_ ;
 wire \i_ibex/id_stage_i/_0318_ ;
 wire \i_ibex/id_stage_i/_0319_ ;
 wire \i_ibex/id_stage_i/_0320_ ;
 wire \i_ibex/id_stage_i/_0321_ ;
 wire \i_ibex/id_stage_i/_0322_ ;
 wire \i_ibex/id_stage_i/_0323_ ;
 wire \i_ibex/id_stage_i/_0324_ ;
 wire \i_ibex/id_stage_i/_0325_ ;
 wire \i_ibex/id_stage_i/_0326_ ;
 wire \i_ibex/id_stage_i/_0327_ ;
 wire \i_ibex/id_stage_i/_0328_ ;
 wire \i_ibex/id_stage_i/_0329_ ;
 wire \i_ibex/id_stage_i/_0330_ ;
 wire \i_ibex/id_stage_i/_0331_ ;
 wire \i_ibex/id_stage_i/_0332_ ;
 wire \i_ibex/id_stage_i/_0333_ ;
 wire net633;
 wire net632;
 wire net631;
 wire net630;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire \i_ibex/id_stage_i/_0342_ ;
 wire \i_ibex/id_stage_i/_0343_ ;
 wire \i_ibex/id_stage_i/_0344_ ;
 wire \i_ibex/id_stage_i/_0345_ ;
 wire \i_ibex/id_stage_i/_0346_ ;
 wire \i_ibex/id_stage_i/_0347_ ;
 wire \i_ibex/id_stage_i/_0348_ ;
 wire net625;
 wire net624;
 wire net623;
 wire net622;
 wire \i_ibex/id_stage_i/_0353_ ;
 wire \i_ibex/id_stage_i/_0354_ ;
 wire \i_ibex/id_stage_i/_0355_ ;
 wire net691;
 wire net690;
 wire net689;
 wire \i_ibex/id_stage_i/_0359_ ;
 wire net688;
 wire \i_ibex/id_stage_i/_0361_ ;
 wire net687;
 wire \i_ibex/id_stage_i/_0363_ ;
 wire \i_ibex/id_stage_i/_0364_ ;
 wire \i_ibex/id_stage_i/_0365_ ;
 wire \i_ibex/id_stage_i/_0366_ ;
 wire net686;
 wire \i_ibex/id_stage_i/_0368_ ;
 wire net685;
 wire net684;
 wire net683;
 wire \i_ibex/id_stage_i/_0372_ ;
 wire \i_ibex/id_stage_i/_0373_ ;
 wire \i_ibex/id_stage_i/_0374_ ;
 wire \i_ibex/id_stage_i/_0375_ ;
 wire \i_ibex/id_stage_i/_0376_ ;
 wire \i_ibex/id_stage_i/_0377_ ;
 wire \i_ibex/id_stage_i/_0378_ ;
 wire \i_ibex/id_stage_i/_0379_ ;
 wire \i_ibex/id_stage_i/_0380_ ;
 wire \i_ibex/id_stage_i/_0381_ ;
 wire \i_ibex/id_stage_i/_0382_ ;
 wire \i_ibex/id_stage_i/_0383_ ;
 wire \i_ibex/id_stage_i/_0384_ ;
 wire \i_ibex/id_stage_i/_0385_ ;
 wire \i_ibex/id_stage_i/_0386_ ;
 wire \i_ibex/id_stage_i/_0387_ ;
 wire \i_ibex/id_stage_i/_0388_ ;
 wire \i_ibex/id_stage_i/_0389_ ;
 wire \i_ibex/id_stage_i/_0390_ ;
 wire \i_ibex/id_stage_i/_0391_ ;
 wire \i_ibex/id_stage_i/_0392_ ;
 wire \i_ibex/id_stage_i/_0393_ ;
 wire \i_ibex/id_stage_i/_0394_ ;
 wire \i_ibex/id_stage_i/_0395_ ;
 wire net682;
 wire \i_ibex/id_stage_i/_0397_ ;
 wire \i_ibex/id_stage_i/_0398_ ;
 wire \i_ibex/id_stage_i/_0399_ ;
 wire \i_ibex/id_stage_i/_0400_ ;
 wire \i_ibex/id_stage_i/_0401_ ;
 wire \i_ibex/id_stage_i/_0402_ ;
 wire \i_ibex/id_stage_i/_0403_ ;
 wire \i_ibex/id_stage_i/_0404_ ;
 wire \i_ibex/id_stage_i/_0405_ ;
 wire \i_ibex/id_stage_i/_0406_ ;
 wire net681;
 wire \i_ibex/id_stage_i/_0408_ ;
 wire \i_ibex/id_stage_i/_0409_ ;
 wire \i_ibex/id_stage_i/_0410_ ;
 wire \i_ibex/id_stage_i/_0411_ ;
 wire net680;
 wire net679;
 wire net678;
 wire \i_ibex/id_stage_i/_0415_ ;
 wire \i_ibex/id_stage_i/_0416_ ;
 wire net677;
 wire net676;
 wire \i_ibex/id_stage_i/_0419_ ;
 wire \i_ibex/id_stage_i/_0420_ ;
 wire \i_ibex/id_stage_i/_0421_ ;
 wire \i_ibex/id_stage_i/_0422_ ;
 wire \i_ibex/id_stage_i/_0423_ ;
 wire \i_ibex/id_stage_i/_0424_ ;
 wire \i_ibex/id_stage_i/_0425_ ;
 wire \i_ibex/id_stage_i/_0426_ ;
 wire \i_ibex/id_stage_i/_0427_ ;
 wire \i_ibex/id_stage_i/_0428_ ;
 wire \i_ibex/id_stage_i/_0429_ ;
 wire \i_ibex/id_stage_i/_0430_ ;
 wire \i_ibex/id_stage_i/_0431_ ;
 wire \i_ibex/id_stage_i/_0432_ ;
 wire \i_ibex/id_stage_i/_0433_ ;
 wire \i_ibex/id_stage_i/_0434_ ;
 wire \i_ibex/id_stage_i/_0435_ ;
 wire \i_ibex/id_stage_i/_0436_ ;
 wire \i_ibex/id_stage_i/_0437_ ;
 wire \i_ibex/id_stage_i/_0438_ ;
 wire \i_ibex/id_stage_i/_0439_ ;
 wire \i_ibex/id_stage_i/_0440_ ;
 wire \i_ibex/id_stage_i/_0441_ ;
 wire \i_ibex/id_stage_i/_0442_ ;
 wire net675;
 wire \i_ibex/id_stage_i/_0444_ ;
 wire \i_ibex/id_stage_i/_0445_ ;
 wire \i_ibex/id_stage_i/_0446_ ;
 wire \i_ibex/id_stage_i/_0447_ ;
 wire \i_ibex/id_stage_i/_0448_ ;
 wire \i_ibex/id_stage_i/_0449_ ;
 wire \i_ibex/id_stage_i/_0450_ ;
 wire \i_ibex/id_stage_i/_0451_ ;
 wire \i_ibex/id_stage_i/_0452_ ;
 wire \i_ibex/id_stage_i/_0453_ ;
 wire net674;
 wire \i_ibex/id_stage_i/_0455_ ;
 wire \i_ibex/id_stage_i/_0456_ ;
 wire \i_ibex/id_stage_i/_0457_ ;
 wire \i_ibex/id_stage_i/_0458_ ;
 wire net673;
 wire net672;
 wire net671;
 wire \i_ibex/id_stage_i/_0462_ ;
 wire \i_ibex/id_stage_i/_0463_ ;
 wire net670;
 wire net669;
 wire \i_ibex/id_stage_i/_0466_ ;
 wire \i_ibex/id_stage_i/_0467_ ;
 wire \i_ibex/id_stage_i/_0468_ ;
 wire \i_ibex/id_stage_i/_0469_ ;
 wire \i_ibex/id_stage_i/_0470_ ;
 wire \i_ibex/id_stage_i/_0471_ ;
 wire \i_ibex/id_stage_i/_0472_ ;
 wire \i_ibex/id_stage_i/_0473_ ;
 wire \i_ibex/id_stage_i/_0474_ ;
 wire \i_ibex/id_stage_i/_0475_ ;
 wire \i_ibex/id_stage_i/_0476_ ;
 wire \i_ibex/id_stage_i/_0477_ ;
 wire \i_ibex/id_stage_i/_0478_ ;
 wire \i_ibex/id_stage_i/_0479_ ;
 wire \i_ibex/id_stage_i/_0480_ ;
 wire \i_ibex/id_stage_i/_0481_ ;
 wire \i_ibex/id_stage_i/_0482_ ;
 wire \i_ibex/id_stage_i/_0483_ ;
 wire \i_ibex/id_stage_i/_0484_ ;
 wire \i_ibex/id_stage_i/_0485_ ;
 wire \i_ibex/id_stage_i/_0486_ ;
 wire \i_ibex/id_stage_i/_0487_ ;
 wire \i_ibex/id_stage_i/_0488_ ;
 wire \i_ibex/id_stage_i/_0489_ ;
 wire \i_ibex/id_stage_i/_0490_ ;
 wire \i_ibex/id_stage_i/_0491_ ;
 wire \i_ibex/id_stage_i/_0492_ ;
 wire \i_ibex/id_stage_i/_0493_ ;
 wire \i_ibex/id_stage_i/_0494_ ;
 wire \i_ibex/id_stage_i/_0495_ ;
 wire \i_ibex/id_stage_i/_0496_ ;
 wire \i_ibex/id_stage_i/_0497_ ;
 wire \i_ibex/id_stage_i/_0498_ ;
 wire \i_ibex/id_stage_i/_0499_ ;
 wire \i_ibex/id_stage_i/_0500_ ;
 wire \i_ibex/id_stage_i/_0501_ ;
 wire \i_ibex/id_stage_i/_0502_ ;
 wire \i_ibex/id_stage_i/_0503_ ;
 wire \i_ibex/id_stage_i/_0504_ ;
 wire \i_ibex/id_stage_i/_0505_ ;
 wire \i_ibex/id_stage_i/_0506_ ;
 wire \i_ibex/id_stage_i/_0507_ ;
 wire \i_ibex/id_stage_i/_0508_ ;
 wire \i_ibex/id_stage_i/_0509_ ;
 wire \i_ibex/id_stage_i/_0510_ ;
 wire \i_ibex/id_stage_i/_0511_ ;
 wire net668;
 wire net667;
 wire \i_ibex/id_stage_i/_0514_ ;
 wire net666;
 wire net665;
 wire \i_ibex/id_stage_i/_0517_ ;
 wire \i_ibex/id_stage_i/_0518_ ;
 wire net664;
 wire \i_ibex/id_stage_i/_0520_ ;
 wire net663;
 wire \i_ibex/id_stage_i/_0522_ ;
 wire \i_ibex/id_stage_i/_0523_ ;
 wire net662;
 wire net661;
 wire net660;
 wire \i_ibex/id_stage_i/_0527_ ;
 wire net659;
 wire \i_ibex/id_stage_i/_0529_ ;
 wire \i_ibex/id_stage_i/_0530_ ;
 wire net658;
 wire \i_ibex/id_stage_i/_0532_ ;
 wire \i_ibex/id_stage_i/_0533_ ;
 wire net657;
 wire net656;
 wire net655;
 wire \i_ibex/id_stage_i/_0537_ ;
 wire net654;
 wire \i_ibex/id_stage_i/_0539_ ;
 wire net653;
 wire \i_ibex/id_stage_i/_0541_ ;
 wire \i_ibex/id_stage_i/_0542_ ;
 wire net652;
 wire \i_ibex/id_stage_i/_0544_ ;
 wire \i_ibex/id_stage_i/_0545_ ;
 wire \i_ibex/id_stage_i/_0546_ ;
 wire \i_ibex/id_stage_i/_0547_ ;
 wire \i_ibex/id_stage_i/_0548_ ;
 wire \i_ibex/id_stage_i/_0549_ ;
 wire \i_ibex/id_stage_i/_0550_ ;
 wire \i_ibex/id_stage_i/_0551_ ;
 wire \i_ibex/id_stage_i/_0552_ ;
 wire \i_ibex/id_stage_i/_0553_ ;
 wire \i_ibex/id_stage_i/_0554_ ;
 wire \i_ibex/id_stage_i/_0555_ ;
 wire \i_ibex/id_stage_i/_0556_ ;
 wire \i_ibex/id_stage_i/_0557_ ;
 wire \i_ibex/id_stage_i/_0558_ ;
 wire \i_ibex/id_stage_i/_0559_ ;
 wire \i_ibex/id_stage_i/_0560_ ;
 wire \i_ibex/id_stage_i/_0561_ ;
 wire \i_ibex/id_stage_i/_0562_ ;
 wire \i_ibex/id_stage_i/_0563_ ;
 wire \i_ibex/id_stage_i/_0564_ ;
 wire \i_ibex/id_stage_i/_0565_ ;
 wire \i_ibex/id_stage_i/_0566_ ;
 wire \i_ibex/id_stage_i/_0567_ ;
 wire \i_ibex/id_stage_i/_0568_ ;
 wire \i_ibex/id_stage_i/_0569_ ;
 wire \i_ibex/id_stage_i/_0570_ ;
 wire \i_ibex/id_stage_i/_0571_ ;
 wire \i_ibex/id_stage_i/_0572_ ;
 wire \i_ibex/id_stage_i/_0573_ ;
 wire \i_ibex/id_stage_i/_0574_ ;
 wire \i_ibex/id_stage_i/_0575_ ;
 wire \i_ibex/id_stage_i/_0576_ ;
 wire \i_ibex/id_stage_i/_0577_ ;
 wire \i_ibex/id_stage_i/_0578_ ;
 wire \i_ibex/id_stage_i/_0579_ ;
 wire \i_ibex/id_stage_i/_0580_ ;
 wire \i_ibex/id_stage_i/_0581_ ;
 wire \i_ibex/id_stage_i/_0582_ ;
 wire \i_ibex/id_stage_i/_0583_ ;
 wire \i_ibex/id_stage_i/_0584_ ;
 wire \i_ibex/id_stage_i/_0585_ ;
 wire \i_ibex/id_stage_i/_0586_ ;
 wire \i_ibex/id_stage_i/_0587_ ;
 wire \i_ibex/id_stage_i/_0588_ ;
 wire \i_ibex/id_stage_i/_0589_ ;
 wire \i_ibex/id_stage_i/_0590_ ;
 wire \i_ibex/id_stage_i/_0591_ ;
 wire \i_ibex/id_stage_i/_0592_ ;
 wire \i_ibex/id_stage_i/_0593_ ;
 wire \i_ibex/id_stage_i/_0594_ ;
 wire \i_ibex/id_stage_i/_0595_ ;
 wire \i_ibex/id_stage_i/_0596_ ;
 wire \i_ibex/id_stage_i/_0597_ ;
 wire \i_ibex/id_stage_i/_0598_ ;
 wire \i_ibex/id_stage_i/_0599_ ;
 wire \i_ibex/id_stage_i/_0600_ ;
 wire \i_ibex/id_stage_i/_0601_ ;
 wire \i_ibex/id_stage_i/_0602_ ;
 wire \i_ibex/id_stage_i/_0603_ ;
 wire \i_ibex/id_stage_i/_0604_ ;
 wire \i_ibex/id_stage_i/_0605_ ;
 wire \i_ibex/id_stage_i/_0606_ ;
 wire \i_ibex/id_stage_i/_0607_ ;
 wire \i_ibex/id_stage_i/_0608_ ;
 wire \i_ibex/id_stage_i/_0609_ ;
 wire \i_ibex/id_stage_i/_0610_ ;
 wire \i_ibex/id_stage_i/_0611_ ;
 wire \i_ibex/id_stage_i/_0612_ ;
 wire \i_ibex/id_stage_i/_0613_ ;
 wire \i_ibex/id_stage_i/_0614_ ;
 wire \i_ibex/id_stage_i/_0615_ ;
 wire \i_ibex/id_stage_i/_0616_ ;
 wire \i_ibex/id_stage_i/_0617_ ;
 wire \i_ibex/id_stage_i/_0618_ ;
 wire \i_ibex/id_stage_i/_0619_ ;
 wire \i_ibex/id_stage_i/_0620_ ;
 wire \i_ibex/id_stage_i/_0621_ ;
 wire \i_ibex/id_stage_i/_0622_ ;
 wire \i_ibex/id_stage_i/_0623_ ;
 wire \i_ibex/id_stage_i/_0624_ ;
 wire \i_ibex/id_stage_i/_0625_ ;
 wire \i_ibex/id_stage_i/_0626_ ;
 wire \i_ibex/id_stage_i/_0627_ ;
 wire \i_ibex/id_stage_i/alu_multicycle_dec ;
 wire \i_ibex/id_stage_i/alu_op_b_mux_sel_dec ;
 wire \i_ibex/id_stage_i/branch_in_dec ;
 wire \i_ibex/id_stage_i/branch_jump_set_done_d ;
 wire \i_ibex/id_stage_i/branch_jump_set_done_q ;
 wire \i_ibex/id_stage_i/branch_set ;
 wire \i_ibex/id_stage_i/branch_set_raw ;
 wire \i_ibex/id_stage_i/branch_set_raw_d ;
 wire \i_ibex/id_stage_i/controller_run ;
 wire \i_ibex/id_stage_i/csr_pipe_flush ;
 wire \i_ibex/id_stage_i/div_en_dec ;
 wire \i_ibex/id_stage_i/dret_insn_dec ;
 wire \i_ibex/id_stage_i/ebrk_insn ;
 wire \i_ibex/id_stage_i/ecall_insn_dec ;
 wire \i_ibex/id_stage_i/flush_id ;
 wire \i_ibex/id_stage_i/id_fsm_q ;
 wire \i_ibex/id_stage_i/illegal_insn_dec ;
 wire \i_ibex/id_stage_i/imm_a_mux_sel ;
 wire \i_ibex/id_stage_i/instr_first_cycle_id_o_$_AND__Y_B ;
 wire \i_ibex/id_stage_i/jump_in_dec ;
 wire \i_ibex/id_stage_i/jump_set ;
 wire \i_ibex/id_stage_i/jump_set_$_AND__Y_B ;
 wire \i_ibex/id_stage_i/jump_set_dec ;
 wire \i_ibex/id_stage_i/lsu_req_dec ;
 wire \i_ibex/id_stage_i/mret_insn_dec ;
 wire \i_ibex/id_stage_i/mult_en_dec ;
 wire \i_ibex/id_stage_i/rf_ren_a_dec ;
 wire \i_ibex/id_stage_i/rf_ren_b_dec ;
 wire \i_ibex/id_stage_i/rf_wdata_sel ;
 wire \i_ibex/id_stage_i/rf_we_dec ;
 wire \i_ibex/id_stage_i/stall_id ;
 wire net380;
 wire \i_ibex/id_stage_i/controller_i/_000_ ;
 wire \i_ibex/id_stage_i/controller_i/_001_ ;
 wire \i_ibex/id_stage_i/controller_i/_002_ ;
 wire \i_ibex/id_stage_i/controller_i/_003_ ;
 wire \i_ibex/id_stage_i/controller_i/_004_ ;
 wire \i_ibex/id_stage_i/controller_i/_005_ ;
 wire \i_ibex/id_stage_i/controller_i/_006_ ;
 wire net621;
 wire \i_ibex/id_stage_i/controller_i/_008_ ;
 wire net620;
 wire net619;
 wire \i_ibex/id_stage_i/controller_i/_011_ ;
 wire \i_ibex/id_stage_i/controller_i/_012_ ;
 wire \i_ibex/id_stage_i/controller_i/_013_ ;
 wire \i_ibex/id_stage_i/controller_i/_014_ ;
 wire \i_ibex/id_stage_i/controller_i/_015_ ;
 wire \i_ibex/id_stage_i/controller_i/_016_ ;
 wire \i_ibex/id_stage_i/controller_i/_017_ ;
 wire \i_ibex/id_stage_i/controller_i/_018_ ;
 wire \i_ibex/id_stage_i/controller_i/_019_ ;
 wire net618;
 wire \i_ibex/id_stage_i/controller_i/_021_ ;
 wire \i_ibex/id_stage_i/controller_i/_022_ ;
 wire \i_ibex/id_stage_i/controller_i/_023_ ;
 wire \i_ibex/id_stage_i/controller_i/_024_ ;
 wire \i_ibex/id_stage_i/controller_i/_025_ ;
 wire \i_ibex/id_stage_i/controller_i/_026_ ;
 wire \i_ibex/id_stage_i/controller_i/_027_ ;
 wire \i_ibex/id_stage_i/controller_i/_028_ ;
 wire net617;
 wire \i_ibex/id_stage_i/controller_i/_030_ ;
 wire \i_ibex/id_stage_i/controller_i/_031_ ;
 wire \i_ibex/id_stage_i/controller_i/_032_ ;
 wire \i_ibex/id_stage_i/controller_i/_033_ ;
 wire \i_ibex/id_stage_i/controller_i/_034_ ;
 wire net616;
 wire \i_ibex/id_stage_i/controller_i/_036_ ;
 wire net615;
 wire \i_ibex/id_stage_i/controller_i/_038_ ;
 wire net614;
 wire \i_ibex/id_stage_i/controller_i/_040_ ;
 wire net613;
 wire \i_ibex/id_stage_i/controller_i/_042_ ;
 wire \i_ibex/id_stage_i/controller_i/_043_ ;
 wire \i_ibex/id_stage_i/controller_i/_044_ ;
 wire \i_ibex/id_stage_i/controller_i/_045_ ;
 wire net612;
 wire net611;
 wire \i_ibex/id_stage_i/controller_i/_048_ ;
 wire \i_ibex/id_stage_i/controller_i/_049_ ;
 wire \i_ibex/id_stage_i/controller_i/_050_ ;
 wire \i_ibex/id_stage_i/controller_i/_051_ ;
 wire \i_ibex/id_stage_i/controller_i/_052_ ;
 wire \i_ibex/id_stage_i/controller_i/_053_ ;
 wire \i_ibex/id_stage_i/controller_i/_054_ ;
 wire \i_ibex/id_stage_i/controller_i/_055_ ;
 wire \i_ibex/id_stage_i/controller_i/_056_ ;
 wire \i_ibex/id_stage_i/controller_i/_057_ ;
 wire \i_ibex/id_stage_i/controller_i/_058_ ;
 wire net610;
 wire \i_ibex/id_stage_i/controller_i/_060_ ;
 wire \i_ibex/id_stage_i/controller_i/_061_ ;
 wire \i_ibex/id_stage_i/controller_i/_062_ ;
 wire \i_ibex/id_stage_i/controller_i/_063_ ;
 wire \i_ibex/id_stage_i/controller_i/_064_ ;
 wire \i_ibex/id_stage_i/controller_i/_065_ ;
 wire \i_ibex/id_stage_i/controller_i/_066_ ;
 wire \i_ibex/id_stage_i/controller_i/_067_ ;
 wire \i_ibex/id_stage_i/controller_i/_068_ ;
 wire \i_ibex/id_stage_i/controller_i/_069_ ;
 wire \i_ibex/id_stage_i/controller_i/_070_ ;
 wire \i_ibex/id_stage_i/controller_i/_071_ ;
 wire \i_ibex/id_stage_i/controller_i/_072_ ;
 wire \i_ibex/id_stage_i/controller_i/_073_ ;
 wire \i_ibex/id_stage_i/controller_i/_074_ ;
 wire \i_ibex/id_stage_i/controller_i/_075_ ;
 wire \i_ibex/id_stage_i/controller_i/_076_ ;
 wire \i_ibex/id_stage_i/controller_i/_077_ ;
 wire \i_ibex/id_stage_i/controller_i/_078_ ;
 wire \i_ibex/id_stage_i/controller_i/_079_ ;
 wire \i_ibex/id_stage_i/controller_i/_080_ ;
 wire net609;
 wire \i_ibex/id_stage_i/controller_i/_082_ ;
 wire \i_ibex/id_stage_i/controller_i/_083_ ;
 wire \i_ibex/id_stage_i/controller_i/_084_ ;
 wire \i_ibex/id_stage_i/controller_i/_085_ ;
 wire \i_ibex/id_stage_i/controller_i/_086_ ;
 wire \i_ibex/id_stage_i/controller_i/_087_ ;
 wire net608;
 wire \i_ibex/id_stage_i/controller_i/_089_ ;
 wire \i_ibex/id_stage_i/controller_i/_090_ ;
 wire \i_ibex/id_stage_i/controller_i/_091_ ;
 wire \i_ibex/id_stage_i/controller_i/_092_ ;
 wire \i_ibex/id_stage_i/controller_i/_093_ ;
 wire net607;
 wire \i_ibex/id_stage_i/controller_i/_095_ ;
 wire \i_ibex/id_stage_i/controller_i/_096_ ;
 wire \i_ibex/id_stage_i/controller_i/_097_ ;
 wire \i_ibex/id_stage_i/controller_i/_098_ ;
 wire \i_ibex/id_stage_i/controller_i/_099_ ;
 wire \i_ibex/id_stage_i/controller_i/_100_ ;
 wire \i_ibex/id_stage_i/controller_i/_101_ ;
 wire \i_ibex/id_stage_i/controller_i/_102_ ;
 wire \i_ibex/id_stage_i/controller_i/_103_ ;
 wire \i_ibex/id_stage_i/controller_i/_104_ ;
 wire \i_ibex/id_stage_i/controller_i/_105_ ;
 wire \i_ibex/id_stage_i/controller_i/_106_ ;
 wire net606;
 wire \i_ibex/id_stage_i/controller_i/_108_ ;
 wire \i_ibex/id_stage_i/controller_i/_109_ ;
 wire \i_ibex/id_stage_i/controller_i/_110_ ;
 wire \i_ibex/id_stage_i/controller_i/_111_ ;
 wire \i_ibex/id_stage_i/controller_i/_112_ ;
 wire \i_ibex/id_stage_i/controller_i/_113_ ;
 wire \i_ibex/id_stage_i/controller_i/_114_ ;
 wire \i_ibex/id_stage_i/controller_i/_115_ ;
 wire \i_ibex/id_stage_i/controller_i/_116_ ;
 wire \i_ibex/id_stage_i/controller_i/_117_ ;
 wire net605;
 wire \i_ibex/id_stage_i/controller_i/_119_ ;
 wire \i_ibex/id_stage_i/controller_i/_120_ ;
 wire \i_ibex/id_stage_i/controller_i/_121_ ;
 wire \i_ibex/id_stage_i/controller_i/_122_ ;
 wire \i_ibex/id_stage_i/controller_i/_123_ ;
 wire \i_ibex/id_stage_i/controller_i/_124_ ;
 wire \i_ibex/id_stage_i/controller_i/_125_ ;
 wire \i_ibex/id_stage_i/controller_i/_126_ ;
 wire \i_ibex/id_stage_i/controller_i/_127_ ;
 wire \i_ibex/id_stage_i/controller_i/_128_ ;
 wire \i_ibex/id_stage_i/controller_i/_129_ ;
 wire \i_ibex/id_stage_i/controller_i/_130_ ;
 wire \i_ibex/id_stage_i/controller_i/_131_ ;
 wire \i_ibex/id_stage_i/controller_i/_132_ ;
 wire \i_ibex/id_stage_i/controller_i/_133_ ;
 wire \i_ibex/id_stage_i/controller_i/_134_ ;
 wire \i_ibex/id_stage_i/controller_i/_135_ ;
 wire net604;
 wire \i_ibex/id_stage_i/controller_i/_137_ ;
 wire \i_ibex/id_stage_i/controller_i/_138_ ;
 wire \i_ibex/id_stage_i/controller_i/_139_ ;
 wire \i_ibex/id_stage_i/controller_i/_140_ ;
 wire \i_ibex/id_stage_i/controller_i/_141_ ;
 wire \i_ibex/id_stage_i/controller_i/_142_ ;
 wire \i_ibex/id_stage_i/controller_i/_143_ ;
 wire \i_ibex/id_stage_i/controller_i/_144_ ;
 wire \i_ibex/id_stage_i/controller_i/_145_ ;
 wire \i_ibex/id_stage_i/controller_i/_146_ ;
 wire \i_ibex/id_stage_i/controller_i/_147_ ;
 wire \i_ibex/id_stage_i/controller_i/_148_ ;
 wire \i_ibex/id_stage_i/controller_i/_149_ ;
 wire \i_ibex/id_stage_i/controller_i/_150_ ;
 wire \i_ibex/id_stage_i/controller_i/_151_ ;
 wire \i_ibex/id_stage_i/controller_i/_152_ ;
 wire \i_ibex/id_stage_i/controller_i/_153_ ;
 wire \i_ibex/id_stage_i/controller_i/_154_ ;
 wire \i_ibex/id_stage_i/controller_i/_155_ ;
 wire \i_ibex/id_stage_i/controller_i/_156_ ;
 wire \i_ibex/id_stage_i/controller_i/_157_ ;
 wire \i_ibex/id_stage_i/controller_i/_158_ ;
 wire \i_ibex/id_stage_i/controller_i/_159_ ;
 wire \i_ibex/id_stage_i/controller_i/_160_ ;
 wire \i_ibex/id_stage_i/controller_i/_161_ ;
 wire \i_ibex/id_stage_i/controller_i/_162_ ;
 wire \i_ibex/id_stage_i/controller_i/_163_ ;
 wire \i_ibex/id_stage_i/controller_i/_164_ ;
 wire \i_ibex/id_stage_i/controller_i/_165_ ;
 wire \i_ibex/id_stage_i/controller_i/_166_ ;
 wire \i_ibex/id_stage_i/controller_i/_167_ ;
 wire \i_ibex/id_stage_i/controller_i/_168_ ;
 wire \i_ibex/id_stage_i/controller_i/_169_ ;
 wire \i_ibex/id_stage_i/controller_i/_170_ ;
 wire \i_ibex/id_stage_i/controller_i/_171_ ;
 wire \i_ibex/id_stage_i/controller_i/_172_ ;
 wire \i_ibex/id_stage_i/controller_i/_173_ ;
 wire \i_ibex/id_stage_i/controller_i/_174_ ;
 wire \i_ibex/id_stage_i/controller_i/_175_ ;
 wire \i_ibex/id_stage_i/controller_i/_176_ ;
 wire \i_ibex/id_stage_i/controller_i/_177_ ;
 wire \i_ibex/id_stage_i/controller_i/_178_ ;
 wire \i_ibex/id_stage_i/controller_i/_179_ ;
 wire \i_ibex/id_stage_i/controller_i/_180_ ;
 wire \i_ibex/id_stage_i/controller_i/_181_ ;
 wire \i_ibex/id_stage_i/controller_i/_182_ ;
 wire \i_ibex/id_stage_i/controller_i/_183_ ;
 wire \i_ibex/id_stage_i/controller_i/_184_ ;
 wire \i_ibex/id_stage_i/controller_i/_185_ ;
 wire \i_ibex/id_stage_i/controller_i/_186_ ;
 wire \i_ibex/id_stage_i/controller_i/_187_ ;
 wire \i_ibex/id_stage_i/controller_i/_188_ ;
 wire \i_ibex/id_stage_i/controller_i/_189_ ;
 wire \i_ibex/id_stage_i/controller_i/_190_ ;
 wire \i_ibex/id_stage_i/controller_i/_191_ ;
 wire \i_ibex/id_stage_i/controller_i/_192_ ;
 wire \i_ibex/id_stage_i/controller_i/_193_ ;
 wire \i_ibex/id_stage_i/controller_i/_194_ ;
 wire \i_ibex/id_stage_i/controller_i/_195_ ;
 wire \i_ibex/id_stage_i/controller_i/_196_ ;
 wire \i_ibex/id_stage_i/controller_i/_197_ ;
 wire \i_ibex/id_stage_i/controller_i/_198_ ;
 wire \i_ibex/id_stage_i/controller_i/_199_ ;
 wire \i_ibex/id_stage_i/controller_i/_200_ ;
 wire \i_ibex/id_stage_i/controller_i/_201_ ;
 wire \i_ibex/id_stage_i/controller_i/_202_ ;
 wire \i_ibex/id_stage_i/controller_i/_203_ ;
 wire \i_ibex/id_stage_i/controller_i/_204_ ;
 wire \i_ibex/id_stage_i/controller_i/_205_ ;
 wire \i_ibex/id_stage_i/controller_i/_206_ ;
 wire \i_ibex/id_stage_i/controller_i/_207_ ;
 wire \i_ibex/id_stage_i/controller_i/_208_ ;
 wire \i_ibex/id_stage_i/controller_i/_209_ ;
 wire \i_ibex/id_stage_i/controller_i/_210_ ;
 wire \i_ibex/id_stage_i/controller_i/_211_ ;
 wire \i_ibex/id_stage_i/controller_i/_212_ ;
 wire \i_ibex/id_stage_i/controller_i/_213_ ;
 wire net603;
 wire \i_ibex/id_stage_i/controller_i/_215_ ;
 wire net602;
 wire \i_ibex/id_stage_i/controller_i/_217_ ;
 wire \i_ibex/id_stage_i/controller_i/_218_ ;
 wire \i_ibex/id_stage_i/controller_i/_219_ ;
 wire net601;
 wire \i_ibex/id_stage_i/controller_i/_221_ ;
 wire \i_ibex/id_stage_i/controller_i/_222_ ;
 wire \i_ibex/id_stage_i/controller_i/_223_ ;
 wire \i_ibex/id_stage_i/controller_i/_224_ ;
 wire \i_ibex/id_stage_i/controller_i/_225_ ;
 wire \i_ibex/id_stage_i/controller_i/_226_ ;
 wire \i_ibex/id_stage_i/controller_i/_227_ ;
 wire \i_ibex/id_stage_i/controller_i/_228_ ;
 wire \i_ibex/id_stage_i/controller_i/_229_ ;
 wire \i_ibex/id_stage_i/controller_i/_230_ ;
 wire \i_ibex/id_stage_i/controller_i/_231_ ;
 wire \i_ibex/id_stage_i/controller_i/_232_ ;
 wire \i_ibex/id_stage_i/controller_i/_233_ ;
 wire \i_ibex/id_stage_i/controller_i/_234_ ;
 wire \i_ibex/id_stage_i/controller_i/_235_ ;
 wire \i_ibex/id_stage_i/controller_i/_236_ ;
 wire \i_ibex/id_stage_i/controller_i/_237_ ;
 wire \i_ibex/id_stage_i/controller_i/_238_ ;
 wire \i_ibex/id_stage_i/controller_i/_239_ ;
 wire \i_ibex/id_stage_i/controller_i/_240_ ;
 wire \i_ibex/id_stage_i/controller_i/_241_ ;
 wire \i_ibex/id_stage_i/controller_i/_242_ ;
 wire \i_ibex/id_stage_i/controller_i/_243_ ;
 wire \i_ibex/id_stage_i/controller_i/_244_ ;
 wire \i_ibex/id_stage_i/controller_i/_245_ ;
 wire \i_ibex/id_stage_i/controller_i/_246_ ;
 wire \i_ibex/id_stage_i/controller_i/_247_ ;
 wire \i_ibex/id_stage_i/controller_i/_248_ ;
 wire \i_ibex/id_stage_i/controller_i/_249_ ;
 wire \i_ibex/id_stage_i/controller_i/_250_ ;
 wire \i_ibex/id_stage_i/controller_i/_251_ ;
 wire \i_ibex/id_stage_i/controller_i/_252_ ;
 wire \i_ibex/id_stage_i/controller_i/_253_ ;
 wire \i_ibex/id_stage_i/controller_i/_254_ ;
 wire \i_ibex/id_stage_i/controller_i/_255_ ;
 wire \i_ibex/id_stage_i/controller_i/_256_ ;
 wire \i_ibex/id_stage_i/controller_i/_257_ ;
 wire \i_ibex/id_stage_i/controller_i/_258_ ;
 wire \i_ibex/id_stage_i/controller_i/_259_ ;
 wire \i_ibex/id_stage_i/controller_i/_260_ ;
 wire \i_ibex/id_stage_i/controller_i/_261_ ;
 wire \i_ibex/id_stage_i/controller_i/_262_ ;
 wire \i_ibex/id_stage_i/controller_i/_263_ ;
 wire \i_ibex/id_stage_i/controller_i/_264_ ;
 wire \i_ibex/id_stage_i/controller_i/_265_ ;
 wire \i_ibex/id_stage_i/controller_i/_266_ ;
 wire \i_ibex/id_stage_i/controller_i/_267_ ;
 wire \i_ibex/id_stage_i/controller_i/_268_ ;
 wire \i_ibex/id_stage_i/controller_i/_269_ ;
 wire \i_ibex/id_stage_i/controller_i/_270_ ;
 wire \i_ibex/id_stage_i/controller_i/_271_ ;
 wire \i_ibex/id_stage_i/controller_i/_272_ ;
 wire \i_ibex/id_stage_i/controller_i/_273_ ;
 wire \i_ibex/id_stage_i/controller_i/_274_ ;
 wire \i_ibex/id_stage_i/controller_i/_275_ ;
 wire \i_ibex/id_stage_i/controller_i/_276_ ;
 wire \i_ibex/id_stage_i/controller_i/_277_ ;
 wire \i_ibex/id_stage_i/controller_i/_278_ ;
 wire \i_ibex/id_stage_i/controller_i/_279_ ;
 wire \i_ibex/id_stage_i/controller_i/_280_ ;
 wire \i_ibex/id_stage_i/controller_i/_281_ ;
 wire \i_ibex/id_stage_i/controller_i/_282_ ;
 wire \i_ibex/id_stage_i/controller_i/_283_ ;
 wire \i_ibex/id_stage_i/controller_i/_284_ ;
 wire \i_ibex/id_stage_i/controller_i/_285_ ;
 wire \i_ibex/id_stage_i/controller_i/_286_ ;
 wire \i_ibex/id_stage_i/controller_i/_287_ ;
 wire \i_ibex/id_stage_i/controller_i/_288_ ;
 wire \i_ibex/id_stage_i/controller_i/_289_ ;
 wire \i_ibex/id_stage_i/controller_i/_290_ ;
 wire \i_ibex/id_stage_i/controller_i/_291_ ;
 wire \i_ibex/id_stage_i/controller_i/_292_ ;
 wire \i_ibex/id_stage_i/controller_i/_293_ ;
 wire \i_ibex/id_stage_i/controller_i/_294_ ;
 wire \i_ibex/id_stage_i/controller_i/_295_ ;
 wire \i_ibex/id_stage_i/controller_i/_296_ ;
 wire \i_ibex/id_stage_i/controller_i/_297_ ;
 wire \i_ibex/id_stage_i/controller_i/_298_ ;
 wire \i_ibex/id_stage_i/controller_i/_299_ ;
 wire \i_ibex/id_stage_i/controller_i/_300_ ;
 wire \i_ibex/id_stage_i/controller_i/_301_ ;
 wire \i_ibex/id_stage_i/controller_i/_302_ ;
 wire \i_ibex/id_stage_i/controller_i/_303_ ;
 wire \i_ibex/id_stage_i/controller_i/_304_ ;
 wire \i_ibex/id_stage_i/controller_i/_305_ ;
 wire \i_ibex/id_stage_i/controller_i/_306_ ;
 wire \i_ibex/id_stage_i/controller_i/_307_ ;
 wire \i_ibex/id_stage_i/controller_i/_308_ ;
 wire \i_ibex/id_stage_i/controller_i/_309_ ;
 wire \i_ibex/id_stage_i/controller_i/_310_ ;
 wire \i_ibex/id_stage_i/controller_i/_311_ ;
 wire \i_ibex/id_stage_i/controller_i/_312_ ;
 wire \i_ibex/id_stage_i/controller_i/_313_ ;
 wire \i_ibex/id_stage_i/controller_i/_314_ ;
 wire \i_ibex/id_stage_i/controller_i/_315_ ;
 wire \i_ibex/id_stage_i/controller_i/_316_ ;
 wire \i_ibex/id_stage_i/controller_i/_317_ ;
 wire \i_ibex/id_stage_i/controller_i/_318_ ;
 wire \i_ibex/id_stage_i/controller_i/_319_ ;
 wire \i_ibex/id_stage_i/controller_i/_320_ ;
 wire \i_ibex/id_stage_i/controller_i/_321_ ;
 wire \i_ibex/id_stage_i/controller_i/_322_ ;
 wire \i_ibex/id_stage_i/controller_i/_323_ ;
 wire \i_ibex/id_stage_i/controller_i/_324_ ;
 wire \i_ibex/id_stage_i/controller_i/_325_ ;
 wire \i_ibex/id_stage_i/controller_i/_326_ ;
 wire \i_ibex/id_stage_i/controller_i/_327_ ;
 wire \i_ibex/id_stage_i/controller_i/_328_ ;
 wire \i_ibex/id_stage_i/controller_i/_329_ ;
 wire \i_ibex/id_stage_i/controller_i/_330_ ;
 wire \i_ibex/id_stage_i/controller_i/_331_ ;
 wire \i_ibex/id_stage_i/controller_i/_332_ ;
 wire \i_ibex/id_stage_i/controller_i/_333_ ;
 wire \i_ibex/id_stage_i/controller_i/_334_ ;
 wire \i_ibex/id_stage_i/controller_i/_335_ ;
 wire \i_ibex/id_stage_i/controller_i/_336_ ;
 wire \i_ibex/id_stage_i/controller_i/_337_ ;
 wire \i_ibex/id_stage_i/controller_i/_338_ ;
 wire \i_ibex/id_stage_i/controller_i/_339_ ;
 wire \i_ibex/id_stage_i/controller_i/_340_ ;
 wire \i_ibex/id_stage_i/controller_i/_341_ ;
 wire \i_ibex/id_stage_i/controller_i/_342_ ;
 wire \i_ibex/id_stage_i/controller_i/_343_ ;
 wire \i_ibex/id_stage_i/controller_i/_344_ ;
 wire \i_ibex/id_stage_i/controller_i/_345_ ;
 wire \i_ibex/id_stage_i/controller_i/_346_ ;
 wire \i_ibex/id_stage_i/controller_i/_347_ ;
 wire \i_ibex/id_stage_i/controller_i/_348_ ;
 wire \i_ibex/id_stage_i/controller_i/_349_ ;
 wire \i_ibex/id_stage_i/controller_i/_350_ ;
 wire \i_ibex/id_stage_i/controller_i/_351_ ;
 wire \i_ibex/id_stage_i/controller_i/_352_ ;
 wire \i_ibex/id_stage_i/controller_i/_353_ ;
 wire \i_ibex/id_stage_i/controller_i/_354_ ;
 wire \i_ibex/id_stage_i/controller_i/_355_ ;
 wire \i_ibex/id_stage_i/controller_i/_356_ ;
 wire \i_ibex/id_stage_i/controller_i/_357_ ;
 wire \i_ibex/id_stage_i/controller_i/_358_ ;
 wire \i_ibex/id_stage_i/controller_i/_359_ ;
 wire \i_ibex/id_stage_i/controller_i/_360_ ;
 wire \i_ibex/id_stage_i/controller_i/_361_ ;
 wire \i_ibex/id_stage_i/controller_i/_362_ ;
 wire \i_ibex/id_stage_i/controller_i/_363_ ;
 wire \i_ibex/id_stage_i/controller_i/_364_ ;
 wire \i_ibex/id_stage_i/controller_i/_365_ ;
 wire \i_ibex/id_stage_i/controller_i/_366_ ;
 wire \i_ibex/id_stage_i/controller_i/_367_ ;
 wire \i_ibex/id_stage_i/controller_i/_368_ ;
 wire \i_ibex/id_stage_i/controller_i/_369_ ;
 wire \i_ibex/id_stage_i/controller_i/_370_ ;
 wire \i_ibex/id_stage_i/controller_i/_371_ ;
 wire \i_ibex/id_stage_i/controller_i/_372_ ;
 wire \i_ibex/id_stage_i/controller_i/_373_ ;
 wire \i_ibex/id_stage_i/controller_i/_374_ ;
 wire \i_ibex/id_stage_i/controller_i/_375_ ;
 wire \i_ibex/id_stage_i/controller_i/_376_ ;
 wire \i_ibex/id_stage_i/controller_i/_377_ ;
 wire \i_ibex/id_stage_i/controller_i/_378_ ;
 wire \i_ibex/id_stage_i/controller_i/_379_ ;
 wire \i_ibex/id_stage_i/controller_i/_380_ ;
 wire \i_ibex/id_stage_i/controller_i/_381_ ;
 wire \i_ibex/id_stage_i/controller_i/_382_ ;
 wire \i_ibex/id_stage_i/controller_i/_383_ ;
 wire \i_ibex/id_stage_i/controller_i/_384_ ;
 wire \i_ibex/id_stage_i/controller_i/_385_ ;
 wire \i_ibex/id_stage_i/controller_i/_386_ ;
 wire \i_ibex/id_stage_i/controller_i/_387_ ;
 wire \i_ibex/id_stage_i/controller_i/_388_ ;
 wire \i_ibex/id_stage_i/controller_i/_389_ ;
 wire \i_ibex/id_stage_i/controller_i/_390_ ;
 wire \i_ibex/id_stage_i/controller_i/_391_ ;
 wire \i_ibex/id_stage_i/controller_i/_392_ ;
 wire \i_ibex/id_stage_i/controller_i/_393_ ;
 wire \i_ibex/id_stage_i/controller_i/_394_ ;
 wire \i_ibex/id_stage_i/controller_i/_395_ ;
 wire \i_ibex/id_stage_i/controller_i/_396_ ;
 wire \i_ibex/id_stage_i/controller_i/_397_ ;
 wire \i_ibex/id_stage_i/controller_i/_398_ ;
 wire \i_ibex/id_stage_i/controller_i/_399_ ;
 wire \i_ibex/id_stage_i/controller_i/_400_ ;
 wire \i_ibex/id_stage_i/controller_i/_401_ ;
 wire \i_ibex/id_stage_i/controller_i/_402_ ;
 wire \i_ibex/id_stage_i/controller_i/_403_ ;
 wire \i_ibex/id_stage_i/controller_i/_404_ ;
 wire \i_ibex/id_stage_i/controller_i/_405_ ;
 wire \i_ibex/id_stage_i/controller_i/_406_ ;
 wire \i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ;
 wire \i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A ;
 wire \i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ;
 wire \i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ;
 wire \i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__B_Y_$_OR__Y_A ;
 wire \i_ibex/id_stage_i/controller_i/do_single_step_d ;
 wire \i_ibex/id_stage_i/controller_i/do_single_step_q ;
 wire \i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_d ;
 wire \i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_q ;
 wire \i_ibex/id_stage_i/controller_i/exc_req_d ;
 wire \i_ibex/id_stage_i/controller_i/exc_req_q ;
 wire \i_ibex/id_stage_i/controller_i/handle_irq_$_AND__Y_A_$_AND__Y_B ;
 wire \i_ibex/id_stage_i/controller_i/illegal_insn_d ;
 wire \i_ibex/id_stage_i/controller_i/illegal_insn_q ;
 wire \i_ibex/id_stage_i/controller_i/load_err_q ;
 wire \i_ibex/id_stage_i/controller_i/store_err_q ;
 wire net595;
 wire \i_ibex/id_stage_i/decoder_i/_001_ ;
 wire \i_ibex/id_stage_i/decoder_i/_002_ ;
 wire \i_ibex/id_stage_i/decoder_i/_003_ ;
 wire net594;
 wire \i_ibex/id_stage_i/decoder_i/_005_ ;
 wire \i_ibex/id_stage_i/decoder_i/_006_ ;
 wire \i_ibex/id_stage_i/decoder_i/_007_ ;
 wire \i_ibex/id_stage_i/decoder_i/_008_ ;
 wire \i_ibex/id_stage_i/decoder_i/_009_ ;
 wire \i_ibex/id_stage_i/decoder_i/_010_ ;
 wire \i_ibex/id_stage_i/decoder_i/_011_ ;
 wire \i_ibex/id_stage_i/decoder_i/_012_ ;
 wire \i_ibex/id_stage_i/decoder_i/_013_ ;
 wire net593;
 wire net592;
 wire \i_ibex/id_stage_i/decoder_i/_016_ ;
 wire \i_ibex/id_stage_i/decoder_i/_017_ ;
 wire \i_ibex/id_stage_i/decoder_i/_018_ ;
 wire \i_ibex/id_stage_i/decoder_i/_019_ ;
 wire net591;
 wire \i_ibex/id_stage_i/decoder_i/_021_ ;
 wire \i_ibex/id_stage_i/decoder_i/_022_ ;
 wire \i_ibex/id_stage_i/decoder_i/_023_ ;
 wire \i_ibex/id_stage_i/decoder_i/_024_ ;
 wire \i_ibex/id_stage_i/decoder_i/_025_ ;
 wire \i_ibex/id_stage_i/decoder_i/_026_ ;
 wire \i_ibex/id_stage_i/decoder_i/_027_ ;
 wire \i_ibex/id_stage_i/decoder_i/_028_ ;
 wire \i_ibex/id_stage_i/decoder_i/_029_ ;
 wire \i_ibex/id_stage_i/decoder_i/_030_ ;
 wire \i_ibex/id_stage_i/decoder_i/_031_ ;
 wire \i_ibex/id_stage_i/decoder_i/_032_ ;
 wire \i_ibex/id_stage_i/decoder_i/_033_ ;
 wire \i_ibex/id_stage_i/decoder_i/_034_ ;
 wire \i_ibex/id_stage_i/decoder_i/_035_ ;
 wire \i_ibex/id_stage_i/decoder_i/_036_ ;
 wire \i_ibex/id_stage_i/decoder_i/_037_ ;
 wire \i_ibex/id_stage_i/decoder_i/_038_ ;
 wire net590;
 wire \i_ibex/id_stage_i/decoder_i/_040_ ;
 wire \i_ibex/id_stage_i/decoder_i/_041_ ;
 wire \i_ibex/id_stage_i/decoder_i/_042_ ;
 wire \i_ibex/id_stage_i/decoder_i/_043_ ;
 wire \i_ibex/id_stage_i/decoder_i/_044_ ;
 wire \i_ibex/id_stage_i/decoder_i/_045_ ;
 wire \i_ibex/id_stage_i/decoder_i/_046_ ;
 wire \i_ibex/id_stage_i/decoder_i/_047_ ;
 wire \i_ibex/id_stage_i/decoder_i/_048_ ;
 wire \i_ibex/id_stage_i/decoder_i/_049_ ;
 wire \i_ibex/id_stage_i/decoder_i/_050_ ;
 wire \i_ibex/id_stage_i/decoder_i/_051_ ;
 wire \i_ibex/id_stage_i/decoder_i/_052_ ;
 wire \i_ibex/id_stage_i/decoder_i/_053_ ;
 wire \i_ibex/id_stage_i/decoder_i/_054_ ;
 wire \i_ibex/id_stage_i/decoder_i/_055_ ;
 wire \i_ibex/id_stage_i/decoder_i/_056_ ;
 wire \i_ibex/id_stage_i/decoder_i/_057_ ;
 wire \i_ibex/id_stage_i/decoder_i/_058_ ;
 wire \i_ibex/id_stage_i/decoder_i/_059_ ;
 wire \i_ibex/id_stage_i/decoder_i/_060_ ;
 wire \i_ibex/id_stage_i/decoder_i/_061_ ;
 wire \i_ibex/id_stage_i/decoder_i/_062_ ;
 wire \i_ibex/id_stage_i/decoder_i/_063_ ;
 wire \i_ibex/id_stage_i/decoder_i/_064_ ;
 wire \i_ibex/id_stage_i/decoder_i/_065_ ;
 wire \i_ibex/id_stage_i/decoder_i/_066_ ;
 wire \i_ibex/id_stage_i/decoder_i/_067_ ;
 wire \i_ibex/id_stage_i/decoder_i/_068_ ;
 wire \i_ibex/id_stage_i/decoder_i/_069_ ;
 wire \i_ibex/id_stage_i/decoder_i/_070_ ;
 wire \i_ibex/id_stage_i/decoder_i/_071_ ;
 wire \i_ibex/id_stage_i/decoder_i/_072_ ;
 wire \i_ibex/id_stage_i/decoder_i/_073_ ;
 wire \i_ibex/id_stage_i/decoder_i/_074_ ;
 wire \i_ibex/id_stage_i/decoder_i/_075_ ;
 wire \i_ibex/id_stage_i/decoder_i/_076_ ;
 wire \i_ibex/id_stage_i/decoder_i/_077_ ;
 wire \i_ibex/id_stage_i/decoder_i/_078_ ;
 wire \i_ibex/id_stage_i/decoder_i/_079_ ;
 wire \i_ibex/id_stage_i/decoder_i/_080_ ;
 wire \i_ibex/id_stage_i/decoder_i/_081_ ;
 wire \i_ibex/id_stage_i/decoder_i/_082_ ;
 wire \i_ibex/id_stage_i/decoder_i/_083_ ;
 wire \i_ibex/id_stage_i/decoder_i/_084_ ;
 wire \i_ibex/id_stage_i/decoder_i/_085_ ;
 wire \i_ibex/id_stage_i/decoder_i/_086_ ;
 wire \i_ibex/id_stage_i/decoder_i/_087_ ;
 wire \i_ibex/id_stage_i/decoder_i/_088_ ;
 wire \i_ibex/id_stage_i/decoder_i/_089_ ;
 wire \i_ibex/id_stage_i/decoder_i/_090_ ;
 wire \i_ibex/id_stage_i/decoder_i/_091_ ;
 wire \i_ibex/id_stage_i/decoder_i/_092_ ;
 wire \i_ibex/id_stage_i/decoder_i/_093_ ;
 wire \i_ibex/id_stage_i/decoder_i/_094_ ;
 wire \i_ibex/id_stage_i/decoder_i/_095_ ;
 wire \i_ibex/id_stage_i/decoder_i/_096_ ;
 wire \i_ibex/id_stage_i/decoder_i/_097_ ;
 wire \i_ibex/id_stage_i/decoder_i/_098_ ;
 wire \i_ibex/id_stage_i/decoder_i/_099_ ;
 wire \i_ibex/id_stage_i/decoder_i/_100_ ;
 wire \i_ibex/id_stage_i/decoder_i/_101_ ;
 wire \i_ibex/id_stage_i/decoder_i/_102_ ;
 wire \i_ibex/id_stage_i/decoder_i/_103_ ;
 wire net589;
 wire \i_ibex/id_stage_i/decoder_i/_105_ ;
 wire \i_ibex/id_stage_i/decoder_i/_106_ ;
 wire net588;
 wire net587;
 wire net586;
 wire \i_ibex/id_stage_i/decoder_i/_110_ ;
 wire \i_ibex/id_stage_i/decoder_i/_111_ ;
 wire \i_ibex/id_stage_i/decoder_i/_112_ ;
 wire \i_ibex/id_stage_i/decoder_i/_113_ ;
 wire \i_ibex/id_stage_i/decoder_i/_114_ ;
 wire \i_ibex/id_stage_i/decoder_i/_115_ ;
 wire net585;
 wire \i_ibex/id_stage_i/decoder_i/_117_ ;
 wire \i_ibex/id_stage_i/decoder_i/_118_ ;
 wire \i_ibex/id_stage_i/decoder_i/_119_ ;
 wire \i_ibex/id_stage_i/decoder_i/_120_ ;
 wire \i_ibex/id_stage_i/decoder_i/_121_ ;
 wire \i_ibex/id_stage_i/decoder_i/_122_ ;
 wire \i_ibex/id_stage_i/decoder_i/_123_ ;
 wire \i_ibex/id_stage_i/decoder_i/_124_ ;
 wire \i_ibex/id_stage_i/decoder_i/_125_ ;
 wire \i_ibex/id_stage_i/decoder_i/_126_ ;
 wire \i_ibex/id_stage_i/decoder_i/_127_ ;
 wire \i_ibex/id_stage_i/decoder_i/_128_ ;
 wire \i_ibex/id_stage_i/decoder_i/_129_ ;
 wire \i_ibex/id_stage_i/decoder_i/_130_ ;
 wire \i_ibex/id_stage_i/decoder_i/_131_ ;
 wire \i_ibex/id_stage_i/decoder_i/_132_ ;
 wire \i_ibex/id_stage_i/decoder_i/_133_ ;
 wire \i_ibex/id_stage_i/decoder_i/_134_ ;
 wire \i_ibex/id_stage_i/decoder_i/_135_ ;
 wire \i_ibex/id_stage_i/decoder_i/_136_ ;
 wire \i_ibex/id_stage_i/decoder_i/_137_ ;
 wire \i_ibex/id_stage_i/decoder_i/_138_ ;
 wire \i_ibex/id_stage_i/decoder_i/_139_ ;
 wire \i_ibex/id_stage_i/decoder_i/_140_ ;
 wire \i_ibex/id_stage_i/decoder_i/_141_ ;
 wire \i_ibex/id_stage_i/decoder_i/_142_ ;
 wire \i_ibex/id_stage_i/decoder_i/_143_ ;
 wire \i_ibex/id_stage_i/decoder_i/_144_ ;
 wire \i_ibex/id_stage_i/decoder_i/_145_ ;
 wire \i_ibex/id_stage_i/decoder_i/_146_ ;
 wire \i_ibex/id_stage_i/decoder_i/_147_ ;
 wire \i_ibex/id_stage_i/decoder_i/_148_ ;
 wire \i_ibex/id_stage_i/decoder_i/_149_ ;
 wire \i_ibex/id_stage_i/decoder_i/_150_ ;
 wire \i_ibex/id_stage_i/decoder_i/_151_ ;
 wire \i_ibex/id_stage_i/decoder_i/_152_ ;
 wire \i_ibex/id_stage_i/decoder_i/_153_ ;
 wire \i_ibex/id_stage_i/decoder_i/_154_ ;
 wire \i_ibex/id_stage_i/decoder_i/_155_ ;
 wire net584;
 wire \i_ibex/id_stage_i/decoder_i/_157_ ;
 wire \i_ibex/id_stage_i/decoder_i/_158_ ;
 wire \i_ibex/id_stage_i/decoder_i/_159_ ;
 wire \i_ibex/id_stage_i/decoder_i/_160_ ;
 wire \i_ibex/id_stage_i/decoder_i/_161_ ;
 wire \i_ibex/id_stage_i/decoder_i/_162_ ;
 wire \i_ibex/id_stage_i/decoder_i/_163_ ;
 wire \i_ibex/id_stage_i/decoder_i/_164_ ;
 wire \i_ibex/id_stage_i/decoder_i/_165_ ;
 wire \i_ibex/id_stage_i/decoder_i/_166_ ;
 wire \i_ibex/id_stage_i/decoder_i/_167_ ;
 wire \i_ibex/id_stage_i/decoder_i/_168_ ;
 wire \i_ibex/id_stage_i/decoder_i/_169_ ;
 wire \i_ibex/id_stage_i/decoder_i/_170_ ;
 wire \i_ibex/id_stage_i/decoder_i/_171_ ;
 wire \i_ibex/id_stage_i/decoder_i/_172_ ;
 wire \i_ibex/id_stage_i/decoder_i/_173_ ;
 wire \i_ibex/id_stage_i/decoder_i/_174_ ;
 wire \i_ibex/id_stage_i/decoder_i/_175_ ;
 wire \i_ibex/id_stage_i/decoder_i/_176_ ;
 wire \i_ibex/id_stage_i/decoder_i/_177_ ;
 wire \i_ibex/id_stage_i/decoder_i/_178_ ;
 wire \i_ibex/id_stage_i/decoder_i/_179_ ;
 wire \i_ibex/id_stage_i/decoder_i/_180_ ;
 wire \i_ibex/id_stage_i/decoder_i/_181_ ;
 wire \i_ibex/id_stage_i/decoder_i/_182_ ;
 wire \i_ibex/id_stage_i/decoder_i/_183_ ;
 wire \i_ibex/id_stage_i/decoder_i/_184_ ;
 wire \i_ibex/id_stage_i/decoder_i/_185_ ;
 wire \i_ibex/id_stage_i/decoder_i/_186_ ;
 wire \i_ibex/id_stage_i/decoder_i/_187_ ;
 wire \i_ibex/id_stage_i/decoder_i/_188_ ;
 wire \i_ibex/id_stage_i/decoder_i/_189_ ;
 wire \i_ibex/id_stage_i/decoder_i/_190_ ;
 wire \i_ibex/id_stage_i/decoder_i/_191_ ;
 wire \i_ibex/id_stage_i/decoder_i/_192_ ;
 wire \i_ibex/id_stage_i/decoder_i/_193_ ;
 wire \i_ibex/id_stage_i/decoder_i/_194_ ;
 wire \i_ibex/id_stage_i/decoder_i/_195_ ;
 wire \i_ibex/id_stage_i/decoder_i/_196_ ;
 wire \i_ibex/id_stage_i/decoder_i/_197_ ;
 wire \i_ibex/id_stage_i/decoder_i/_198_ ;
 wire \i_ibex/id_stage_i/decoder_i/_199_ ;
 wire \i_ibex/id_stage_i/decoder_i/_200_ ;
 wire \i_ibex/id_stage_i/decoder_i/_201_ ;
 wire \i_ibex/id_stage_i/decoder_i/_202_ ;
 wire \i_ibex/id_stage_i/decoder_i/_203_ ;
 wire \i_ibex/id_stage_i/decoder_i/_204_ ;
 wire \i_ibex/id_stage_i/decoder_i/_205_ ;
 wire \i_ibex/id_stage_i/decoder_i/_206_ ;
 wire \i_ibex/id_stage_i/decoder_i/_207_ ;
 wire \i_ibex/id_stage_i/decoder_i/_208_ ;
 wire \i_ibex/id_stage_i/decoder_i/_209_ ;
 wire \i_ibex/id_stage_i/decoder_i/_210_ ;
 wire \i_ibex/id_stage_i/decoder_i/_211_ ;
 wire \i_ibex/id_stage_i/decoder_i/_212_ ;
 wire \i_ibex/id_stage_i/decoder_i/_213_ ;
 wire \i_ibex/id_stage_i/decoder_i/_214_ ;
 wire \i_ibex/id_stage_i/decoder_i/_215_ ;
 wire \i_ibex/id_stage_i/decoder_i/_216_ ;
 wire \i_ibex/id_stage_i/decoder_i/_217_ ;
 wire \i_ibex/id_stage_i/decoder_i/_218_ ;
 wire \i_ibex/id_stage_i/decoder_i/_219_ ;
 wire \i_ibex/id_stage_i/decoder_i/_220_ ;
 wire \i_ibex/id_stage_i/decoder_i/_221_ ;
 wire \i_ibex/id_stage_i/decoder_i/_222_ ;
 wire \i_ibex/id_stage_i/decoder_i/_223_ ;
 wire \i_ibex/id_stage_i/decoder_i/_224_ ;
 wire \i_ibex/id_stage_i/decoder_i/_225_ ;
 wire \i_ibex/id_stage_i/decoder_i/_226_ ;
 wire \i_ibex/id_stage_i/decoder_i/_227_ ;
 wire net600;
 wire net599;
 wire net598;
 wire net597;
 wire net596;
 wire \i_ibex/id_stage_i/decoder_i/_233_ ;
 wire \i_ibex/id_stage_i/decoder_i/_234_ ;
 wire \i_ibex/id_stage_i/decoder_i/_235_ ;
 wire \i_ibex/id_stage_i/decoder_i/_236_ ;
 wire \i_ibex/if_stage_i/_000_ ;
 wire \i_ibex/if_stage_i/_001_ ;
 wire \i_ibex/if_stage_i/_002_ ;
 wire \i_ibex/if_stage_i/_003_ ;
 wire \i_ibex/if_stage_i/_004_ ;
 wire \i_ibex/if_stage_i/_005_ ;
 wire \i_ibex/if_stage_i/_006_ ;
 wire \i_ibex/if_stage_i/_007_ ;
 wire \i_ibex/if_stage_i/_008_ ;
 wire \i_ibex/if_stage_i/_009_ ;
 wire \i_ibex/if_stage_i/_010_ ;
 wire \i_ibex/if_stage_i/_011_ ;
 wire \i_ibex/if_stage_i/_012_ ;
 wire \i_ibex/if_stage_i/_013_ ;
 wire \i_ibex/if_stage_i/_014_ ;
 wire \i_ibex/if_stage_i/_015_ ;
 wire \i_ibex/if_stage_i/_016_ ;
 wire \i_ibex/if_stage_i/_017_ ;
 wire \i_ibex/if_stage_i/_018_ ;
 wire \i_ibex/if_stage_i/_019_ ;
 wire \i_ibex/if_stage_i/_020_ ;
 wire \i_ibex/if_stage_i/_021_ ;
 wire \i_ibex/if_stage_i/_022_ ;
 wire \i_ibex/if_stage_i/_023_ ;
 wire \i_ibex/if_stage_i/_024_ ;
 wire \i_ibex/if_stage_i/_025_ ;
 wire \i_ibex/if_stage_i/_026_ ;
 wire \i_ibex/if_stage_i/_027_ ;
 wire \i_ibex/if_stage_i/_028_ ;
 wire \i_ibex/if_stage_i/_029_ ;
 wire \i_ibex/if_stage_i/_030_ ;
 wire \i_ibex/if_stage_i/_031_ ;
 wire \i_ibex/if_stage_i/_032_ ;
 wire \i_ibex/if_stage_i/_033_ ;
 wire \i_ibex/if_stage_i/_034_ ;
 wire \i_ibex/if_stage_i/_035_ ;
 wire \i_ibex/if_stage_i/_036_ ;
 wire \i_ibex/if_stage_i/_037_ ;
 wire \i_ibex/if_stage_i/_038_ ;
 wire \i_ibex/if_stage_i/_039_ ;
 wire \i_ibex/if_stage_i/_040_ ;
 wire \i_ibex/if_stage_i/_041_ ;
 wire \i_ibex/if_stage_i/_042_ ;
 wire \i_ibex/if_stage_i/_043_ ;
 wire \i_ibex/if_stage_i/_044_ ;
 wire \i_ibex/if_stage_i/_045_ ;
 wire \i_ibex/if_stage_i/_046_ ;
 wire \i_ibex/if_stage_i/_047_ ;
 wire \i_ibex/if_stage_i/_048_ ;
 wire \i_ibex/if_stage_i/_049_ ;
 wire \i_ibex/if_stage_i/_050_ ;
 wire \i_ibex/if_stage_i/_051_ ;
 wire \i_ibex/if_stage_i/_052_ ;
 wire \i_ibex/if_stage_i/_053_ ;
 wire \i_ibex/if_stage_i/_054_ ;
 wire \i_ibex/if_stage_i/_055_ ;
 wire \i_ibex/if_stage_i/_056_ ;
 wire \i_ibex/if_stage_i/_057_ ;
 wire \i_ibex/if_stage_i/_058_ ;
 wire \i_ibex/if_stage_i/_059_ ;
 wire \i_ibex/if_stage_i/_060_ ;
 wire \i_ibex/if_stage_i/_061_ ;
 wire \i_ibex/if_stage_i/_062_ ;
 wire \i_ibex/if_stage_i/_063_ ;
 wire \i_ibex/if_stage_i/_064_ ;
 wire \i_ibex/if_stage_i/_065_ ;
 wire \i_ibex/if_stage_i/_066_ ;
 wire \i_ibex/if_stage_i/_067_ ;
 wire \i_ibex/if_stage_i/_068_ ;
 wire \i_ibex/if_stage_i/_069_ ;
 wire \i_ibex/if_stage_i/_070_ ;
 wire \i_ibex/if_stage_i/_071_ ;
 wire \i_ibex/if_stage_i/_072_ ;
 wire \i_ibex/if_stage_i/_073_ ;
 wire \i_ibex/if_stage_i/_074_ ;
 wire \i_ibex/if_stage_i/_075_ ;
 wire \i_ibex/if_stage_i/_076_ ;
 wire \i_ibex/if_stage_i/_077_ ;
 wire \i_ibex/if_stage_i/_078_ ;
 wire \i_ibex/if_stage_i/_079_ ;
 wire \i_ibex/if_stage_i/_080_ ;
 wire \i_ibex/if_stage_i/_081_ ;
 wire \i_ibex/if_stage_i/_082_ ;
 wire \i_ibex/if_stage_i/_083_ ;
 wire \i_ibex/if_stage_i/_084_ ;
 wire net583;
 wire net582;
 wire net581;
 wire net580;
 wire net579;
 wire net578;
 wire \i_ibex/if_stage_i/_091_ ;
 wire \i_ibex/if_stage_i/_092_ ;
 wire \i_ibex/if_stage_i/_093_ ;
 wire net577;
 wire net576;
 wire \i_ibex/if_stage_i/_096_ ;
 wire net575;
 wire \i_ibex/if_stage_i/_098_ ;
 wire net574;
 wire \i_ibex/if_stage_i/_100_ ;
 wire net573;
 wire \i_ibex/if_stage_i/_102_ ;
 wire net572;
 wire \i_ibex/if_stage_i/_104_ ;
 wire \i_ibex/if_stage_i/_105_ ;
 wire \i_ibex/if_stage_i/_106_ ;
 wire \i_ibex/if_stage_i/_107_ ;
 wire net571;
 wire net570;
 wire \i_ibex/if_stage_i/_110_ ;
 wire \i_ibex/if_stage_i/_111_ ;
 wire \i_ibex/if_stage_i/_112_ ;
 wire net569;
 wire \i_ibex/if_stage_i/_114_ ;
 wire \i_ibex/if_stage_i/_115_ ;
 wire \i_ibex/if_stage_i/_116_ ;
 wire \i_ibex/if_stage_i/_117_ ;
 wire \i_ibex/if_stage_i/_118_ ;
 wire \i_ibex/if_stage_i/_119_ ;
 wire \i_ibex/if_stage_i/_120_ ;
 wire net568;
 wire \i_ibex/if_stage_i/_122_ ;
 wire net567;
 wire \i_ibex/if_stage_i/_124_ ;
 wire \i_ibex/if_stage_i/_125_ ;
 wire \i_ibex/if_stage_i/_126_ ;
 wire \i_ibex/if_stage_i/_127_ ;
 wire \i_ibex/if_stage_i/_128_ ;
 wire \i_ibex/if_stage_i/_129_ ;
 wire \i_ibex/if_stage_i/_130_ ;
 wire \i_ibex/if_stage_i/_131_ ;
 wire \i_ibex/if_stage_i/_132_ ;
 wire \i_ibex/if_stage_i/_133_ ;
 wire \i_ibex/if_stage_i/_134_ ;
 wire \i_ibex/if_stage_i/_135_ ;
 wire \i_ibex/if_stage_i/_136_ ;
 wire \i_ibex/if_stage_i/_137_ ;
 wire \i_ibex/if_stage_i/_138_ ;
 wire \i_ibex/if_stage_i/_139_ ;
 wire \i_ibex/if_stage_i/_140_ ;
 wire \i_ibex/if_stage_i/_141_ ;
 wire \i_ibex/if_stage_i/_142_ ;
 wire \i_ibex/if_stage_i/_143_ ;
 wire \i_ibex/if_stage_i/_144_ ;
 wire \i_ibex/if_stage_i/_145_ ;
 wire \i_ibex/if_stage_i/_146_ ;
 wire \i_ibex/if_stage_i/_147_ ;
 wire \i_ibex/if_stage_i/_148_ ;
 wire \i_ibex/if_stage_i/_149_ ;
 wire net566;
 wire \i_ibex/if_stage_i/_151_ ;
 wire \i_ibex/if_stage_i/_152_ ;
 wire net565;
 wire \i_ibex/if_stage_i/_154_ ;
 wire \i_ibex/if_stage_i/_155_ ;
 wire \i_ibex/if_stage_i/_156_ ;
 wire \i_ibex/if_stage_i/_157_ ;
 wire \i_ibex/if_stage_i/_158_ ;
 wire \i_ibex/if_stage_i/_159_ ;
 wire \i_ibex/if_stage_i/_160_ ;
 wire net564;
 wire \i_ibex/if_stage_i/_162_ ;
 wire \i_ibex/if_stage_i/_163_ ;
 wire \i_ibex/if_stage_i/_164_ ;
 wire \i_ibex/if_stage_i/_165_ ;
 wire \i_ibex/if_stage_i/_166_ ;
 wire \i_ibex/if_stage_i/_167_ ;
 wire \i_ibex/if_stage_i/_168_ ;
 wire \i_ibex/if_stage_i/_169_ ;
 wire \i_ibex/if_stage_i/_170_ ;
 wire \i_ibex/if_stage_i/_171_ ;
 wire \i_ibex/if_stage_i/_172_ ;
 wire \i_ibex/if_stage_i/_173_ ;
 wire \i_ibex/if_stage_i/_174_ ;
 wire \i_ibex/if_stage_i/_175_ ;
 wire \i_ibex/if_stage_i/_176_ ;
 wire \i_ibex/if_stage_i/_177_ ;
 wire \i_ibex/if_stage_i/_178_ ;
 wire \i_ibex/if_stage_i/_179_ ;
 wire \i_ibex/if_stage_i/_180_ ;
 wire \i_ibex/if_stage_i/_181_ ;
 wire \i_ibex/if_stage_i/_182_ ;
 wire \i_ibex/if_stage_i/_183_ ;
 wire \i_ibex/if_stage_i/_184_ ;
 wire \i_ibex/if_stage_i/_185_ ;
 wire \i_ibex/if_stage_i/_186_ ;
 wire \i_ibex/if_stage_i/_187_ ;
 wire \i_ibex/if_stage_i/_188_ ;
 wire \i_ibex/if_stage_i/_189_ ;
 wire \i_ibex/if_stage_i/_190_ ;
 wire \i_ibex/if_stage_i/_191_ ;
 wire \i_ibex/if_stage_i/_192_ ;
 wire net563;
 wire net562;
 wire net561;
 wire \i_ibex/if_stage_i/_196_ ;
 wire \i_ibex/if_stage_i/_197_ ;
 wire \i_ibex/if_stage_i/_198_ ;
 wire \i_ibex/if_stage_i/_199_ ;
 wire net560;
 wire \i_ibex/if_stage_i/_201_ ;
 wire net559;
 wire \i_ibex/if_stage_i/_203_ ;
 wire \i_ibex/if_stage_i/_204_ ;
 wire \i_ibex/if_stage_i/_205_ ;
 wire \i_ibex/if_stage_i/_206_ ;
 wire \i_ibex/if_stage_i/_207_ ;
 wire \i_ibex/if_stage_i/_208_ ;
 wire \i_ibex/if_stage_i/_209_ ;
 wire \i_ibex/if_stage_i/_210_ ;
 wire net558;
 wire \i_ibex/if_stage_i/_212_ ;
 wire net557;
 wire \i_ibex/if_stage_i/_214_ ;
 wire \i_ibex/if_stage_i/_215_ ;
 wire \i_ibex/if_stage_i/_216_ ;
 wire \i_ibex/if_stage_i/_217_ ;
 wire \i_ibex/if_stage_i/_218_ ;
 wire \i_ibex/if_stage_i/_219_ ;
 wire \i_ibex/if_stage_i/_220_ ;
 wire \i_ibex/if_stage_i/_221_ ;
 wire \i_ibex/if_stage_i/_222_ ;
 wire \i_ibex/if_stage_i/_223_ ;
 wire \i_ibex/if_stage_i/_224_ ;
 wire \i_ibex/if_stage_i/_225_ ;
 wire \i_ibex/if_stage_i/_226_ ;
 wire \i_ibex/if_stage_i/_227_ ;
 wire \i_ibex/if_stage_i/_228_ ;
 wire \i_ibex/if_stage_i/_229_ ;
 wire \i_ibex/if_stage_i/_230_ ;
 wire \i_ibex/if_stage_i/_231_ ;
 wire \i_ibex/if_stage_i/_232_ ;
 wire \i_ibex/if_stage_i/_233_ ;
 wire \i_ibex/if_stage_i/_234_ ;
 wire \i_ibex/if_stage_i/_235_ ;
 wire \i_ibex/if_stage_i/_236_ ;
 wire \i_ibex/if_stage_i/_237_ ;
 wire \i_ibex/if_stage_i/_238_ ;
 wire \i_ibex/if_stage_i/_239_ ;
 wire \i_ibex/if_stage_i/_240_ ;
 wire \i_ibex/if_stage_i/_241_ ;
 wire \i_ibex/if_stage_i/_242_ ;
 wire \i_ibex/if_stage_i/_243_ ;
 wire \i_ibex/if_stage_i/_244_ ;
 wire \i_ibex/if_stage_i/_245_ ;
 wire \i_ibex/if_stage_i/_246_ ;
 wire \i_ibex/if_stage_i/_247_ ;
 wire \i_ibex/if_stage_i/_248_ ;
 wire \i_ibex/if_stage_i/_249_ ;
 wire \i_ibex/if_stage_i/_250_ ;
 wire net556;
 wire \i_ibex/if_stage_i/_252_ ;
 wire \i_ibex/if_stage_i/_253_ ;
 wire \i_ibex/if_stage_i/_254_ ;
 wire \i_ibex/if_stage_i/_255_ ;
 wire \i_ibex/if_stage_i/_256_ ;
 wire \i_ibex/if_stage_i/_257_ ;
 wire \i_ibex/if_stage_i/_258_ ;
 wire \i_ibex/if_stage_i/_259_ ;
 wire \i_ibex/if_stage_i/_260_ ;
 wire \i_ibex/if_stage_i/_261_ ;
 wire \i_ibex/if_stage_i/_262_ ;
 wire \i_ibex/if_stage_i/_263_ ;
 wire \i_ibex/if_stage_i/_264_ ;
 wire \i_ibex/if_stage_i/_265_ ;
 wire \i_ibex/if_stage_i/_266_ ;
 wire \i_ibex/if_stage_i/_267_ ;
 wire \i_ibex/if_stage_i/_268_ ;
 wire \i_ibex/if_stage_i/_269_ ;
 wire \i_ibex/if_stage_i/_270_ ;
 wire \i_ibex/if_stage_i/_271_ ;
 wire \i_ibex/if_stage_i/_272_ ;
 wire \i_ibex/if_stage_i/_273_ ;
 wire \i_ibex/if_stage_i/_274_ ;
 wire \i_ibex/if_stage_i/_275_ ;
 wire \i_ibex/if_stage_i/_276_ ;
 wire \i_ibex/if_stage_i/_277_ ;
 wire \i_ibex/if_stage_i/_278_ ;
 wire \i_ibex/if_stage_i/_279_ ;
 wire \i_ibex/if_stage_i/_280_ ;
 wire \i_ibex/if_stage_i/_281_ ;
 wire \i_ibex/if_stage_i/_282_ ;
 wire \i_ibex/if_stage_i/_283_ ;
 wire \i_ibex/if_stage_i/_284_ ;
 wire \i_ibex/if_stage_i/_285_ ;
 wire \i_ibex/if_stage_i/_286_ ;
 wire \i_ibex/if_stage_i/_287_ ;
 wire \i_ibex/if_stage_i/_288_ ;
 wire \i_ibex/if_stage_i/_289_ ;
 wire \i_ibex/if_stage_i/_290_ ;
 wire \i_ibex/if_stage_i/_291_ ;
 wire \i_ibex/if_stage_i/_292_ ;
 wire \i_ibex/if_stage_i/_293_ ;
 wire \i_ibex/if_stage_i/_294_ ;
 wire \i_ibex/if_stage_i/_295_ ;
 wire \i_ibex/if_stage_i/_296_ ;
 wire \i_ibex/if_stage_i/_297_ ;
 wire \i_ibex/if_stage_i/_298_ ;
 wire \i_ibex/if_stage_i/_299_ ;
 wire \i_ibex/if_stage_i/_300_ ;
 wire \i_ibex/if_stage_i/_301_ ;
 wire \i_ibex/if_stage_i/_302_ ;
 wire \i_ibex/if_stage_i/_303_ ;
 wire \i_ibex/if_stage_i/_304_ ;
 wire \i_ibex/if_stage_i/_305_ ;
 wire \i_ibex/if_stage_i/_306_ ;
 wire \i_ibex/if_stage_i/_307_ ;
 wire \i_ibex/if_stage_i/_308_ ;
 wire \i_ibex/if_stage_i/_309_ ;
 wire \i_ibex/if_stage_i/_310_ ;
 wire \i_ibex/if_stage_i/_311_ ;
 wire \i_ibex/if_stage_i/_312_ ;
 wire \i_ibex/if_stage_i/_313_ ;
 wire \i_ibex/if_stage_i/_314_ ;
 wire \i_ibex/if_stage_i/_315_ ;
 wire \i_ibex/if_stage_i/_316_ ;
 wire \i_ibex/if_stage_i/_317_ ;
 wire \i_ibex/if_stage_i/_318_ ;
 wire \i_ibex/if_stage_i/_319_ ;
 wire \i_ibex/if_stage_i/_320_ ;
 wire \i_ibex/if_stage_i/_321_ ;
 wire \i_ibex/if_stage_i/_322_ ;
 wire \i_ibex/if_stage_i/_323_ ;
 wire \i_ibex/if_stage_i/_324_ ;
 wire \i_ibex/if_stage_i/_325_ ;
 wire \i_ibex/if_stage_i/_326_ ;
 wire \i_ibex/if_stage_i/_327_ ;
 wire \i_ibex/if_stage_i/_328_ ;
 wire \i_ibex/if_stage_i/_329_ ;
 wire \i_ibex/if_stage_i/_330_ ;
 wire \i_ibex/if_stage_i/_331_ ;
 wire \i_ibex/if_stage_i/_332_ ;
 wire \i_ibex/if_stage_i/_333_ ;
 wire \i_ibex/if_stage_i/_334_ ;
 wire \i_ibex/if_stage_i/_335_ ;
 wire \i_ibex/if_stage_i/_336_ ;
 wire \i_ibex/if_stage_i/_337_ ;
 wire \i_ibex/if_stage_i/_338_ ;
 wire \i_ibex/if_stage_i/_339_ ;
 wire \i_ibex/if_stage_i/_340_ ;
 wire net555;
 wire \i_ibex/if_stage_i/_342_ ;
 wire \i_ibex/if_stage_i/_343_ ;
 wire \i_ibex/if_stage_i/_344_ ;
 wire \i_ibex/if_stage_i/_345_ ;
 wire \i_ibex/if_stage_i/_346_ ;
 wire net553;
 wire net552;
 wire net551;
 wire net550;
 wire net549;
 wire \i_ibex/if_stage_i/_352_ ;
 wire net548;
 wire net547;
 wire \i_ibex/if_stage_i/_355_ ;
 wire \i_ibex/if_stage_i/_356_ ;
 wire \i_ibex/if_stage_i/_357_ ;
 wire \i_ibex/if_stage_i/_358_ ;
 wire \i_ibex/if_stage_i/_359_ ;
 wire \i_ibex/if_stage_i/_360_ ;
 wire \i_ibex/if_stage_i/_361_ ;
 wire \i_ibex/if_stage_i/_362_ ;
 wire \i_ibex/if_stage_i/_363_ ;
 wire \i_ibex/if_stage_i/_364_ ;
 wire \i_ibex/if_stage_i/_365_ ;
 wire \i_ibex/if_stage_i/_366_ ;
 wire \i_ibex/if_stage_i/_367_ ;
 wire \i_ibex/if_stage_i/_368_ ;
 wire \i_ibex/if_stage_i/_369_ ;
 wire \i_ibex/if_stage_i/_370_ ;
 wire \i_ibex/if_stage_i/_371_ ;
 wire \i_ibex/if_stage_i/_372_ ;
 wire \i_ibex/if_stage_i/_373_ ;
 wire \i_ibex/if_stage_i/_374_ ;
 wire \i_ibex/if_stage_i/_375_ ;
 wire \i_ibex/if_stage_i/_376_ ;
 wire \i_ibex/if_stage_i/_377_ ;
 wire \i_ibex/if_stage_i/_378_ ;
 wire \i_ibex/if_stage_i/_379_ ;
 wire \i_ibex/if_stage_i/_380_ ;
 wire \i_ibex/if_stage_i/_381_ ;
 wire \i_ibex/if_stage_i/_382_ ;
 wire \i_ibex/if_stage_i/_383_ ;
 wire \i_ibex/if_stage_i/_384_ ;
 wire \i_ibex/if_stage_i/_385_ ;
 wire \i_ibex/if_stage_i/_386_ ;
 wire \i_ibex/if_stage_i/_387_ ;
 wire \i_ibex/if_stage_i/_388_ ;
 wire \i_ibex/if_stage_i/_389_ ;
 wire \i_ibex/if_stage_i/_390_ ;
 wire \i_ibex/if_stage_i/_391_ ;
 wire \i_ibex/if_stage_i/_392_ ;
 wire \i_ibex/if_stage_i/_393_ ;
 wire \i_ibex/if_stage_i/_394_ ;
 wire \i_ibex/if_stage_i/_395_ ;
 wire \i_ibex/if_stage_i/_396_ ;
 wire \i_ibex/if_stage_i/_397_ ;
 wire \i_ibex/if_stage_i/_398_ ;
 wire \i_ibex/if_stage_i/_399_ ;
 wire \i_ibex/if_stage_i/_400_ ;
 wire \i_ibex/if_stage_i/_401_ ;
 wire \i_ibex/if_stage_i/_402_ ;
 wire \i_ibex/if_stage_i/_403_ ;
 wire \i_ibex/if_stage_i/_404_ ;
 wire \i_ibex/if_stage_i/_405_ ;
 wire \i_ibex/if_stage_i/_406_ ;
 wire \i_ibex/if_stage_i/_407_ ;
 wire \i_ibex/if_stage_i/_408_ ;
 wire \i_ibex/if_stage_i/_409_ ;
 wire \i_ibex/if_stage_i/_410_ ;
 wire \i_ibex/if_stage_i/_411_ ;
 wire \i_ibex/if_stage_i/_412_ ;
 wire \i_ibex/if_stage_i/_413_ ;
 wire \i_ibex/if_stage_i/_414_ ;
 wire \i_ibex/if_stage_i/_415_ ;
 wire \i_ibex/if_stage_i/_416_ ;
 wire \i_ibex/if_stage_i/_417_ ;
 wire \i_ibex/if_stage_i/_418_ ;
 wire \i_ibex/if_stage_i/_419_ ;
 wire \i_ibex/if_stage_i/_420_ ;
 wire \i_ibex/if_stage_i/_421_ ;
 wire \i_ibex/if_stage_i/_422_ ;
 wire \i_ibex/if_stage_i/_423_ ;
 wire \i_ibex/if_stage_i/_424_ ;
 wire \i_ibex/if_stage_i/_425_ ;
 wire \i_ibex/if_stage_i/_426_ ;
 wire \i_ibex/if_stage_i/_427_ ;
 wire \i_ibex/if_stage_i/_428_ ;
 wire \i_ibex/if_stage_i/_429_ ;
 wire \i_ibex/if_stage_i/_430_ ;
 wire \i_ibex/if_stage_i/_431_ ;
 wire \i_ibex/if_stage_i/_432_ ;
 wire \i_ibex/if_stage_i/_433_ ;
 wire \i_ibex/if_stage_i/_434_ ;
 wire \i_ibex/if_stage_i/_435_ ;
 wire \i_ibex/if_stage_i/_436_ ;
 wire \i_ibex/if_stage_i/_437_ ;
 wire \i_ibex/if_stage_i/_438_ ;
 wire \i_ibex/if_stage_i/_439_ ;
 wire \i_ibex/if_stage_i/_440_ ;
 wire net379;
 wire \i_ibex/if_stage_i/compressed_decoder_i_valid_i ;
 wire \i_ibex/if_stage_i/fetch_err ;
 wire \i_ibex/if_stage_i/fetch_err_plus2 ;
 wire \i_ibex/if_stage_i/fetch_valid ;
 wire net554;
 wire \i_ibex/if_stage_i/illegal_c_insn ;
 wire \i_ibex/if_stage_i/instr_is_compressed ;
 wire \i_ibex/if_stage_i/instr_valid_id_d ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_000_ ;
 wire net529;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_002_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_003_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_004_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_005_ ;
 wire net528;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_007_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_008_ ;
 wire net527;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_010_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_011_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_012_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_013_ ;
 wire net526;
 wire net525;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_016_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_017_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_018_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_019_ ;
 wire net524;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_021_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_022_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_023_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_024_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_025_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_026_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_027_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_028_ ;
 wire net523;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_030_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_031_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_032_ ;
 wire net522;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_034_ ;
 wire net521;
 wire net520;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_037_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_038_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_039_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_040_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_041_ ;
 wire net519;
 wire net518;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_044_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_045_ ;
 wire net517;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_047_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_048_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_049_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_050_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_051_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_052_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_053_ ;
 wire net516;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_055_ ;
 wire net515;
 wire net514;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_058_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_059_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_060_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_061_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_062_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_063_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_064_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_065_ ;
 wire net513;
 wire net512;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_068_ ;
 wire net511;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_070_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_071_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_072_ ;
 wire net510;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_074_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_075_ ;
 wire net509;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_077_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_078_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_079_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_080_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_081_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_082_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_083_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_084_ ;
 wire net508;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_086_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_087_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_088_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_089_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_090_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_091_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_092_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_093_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_094_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_095_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_096_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_097_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_098_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_099_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_100_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_101_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_102_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_103_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_104_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_105_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_106_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_107_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_108_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_109_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_110_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_111_ ;
 wire net507;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_113_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_114_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_115_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_116_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_117_ ;
 wire net506;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_119_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_120_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_121_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_122_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_123_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_124_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_125_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_126_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_127_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_128_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_129_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_130_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_131_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_132_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_133_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_134_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_135_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_136_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_137_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_138_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_139_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_140_ ;
 wire net505;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_142_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_143_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_144_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_145_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_146_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_147_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_148_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_149_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_150_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_151_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_152_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_153_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_154_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_155_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_156_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_157_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_158_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_159_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_160_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_161_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_162_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_163_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_164_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_165_ ;
 wire net504;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_167_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_168_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_169_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_170_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_171_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_172_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_173_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_174_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_175_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_176_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_177_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_178_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_179_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_180_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_181_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_182_ ;
 wire net503;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_184_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_185_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_186_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_187_ ;
 wire net502;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_189_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_190_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_191_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_192_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_193_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_194_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_195_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_196_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_197_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_198_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_199_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_200_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_201_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_202_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_203_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_204_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_205_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_206_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_207_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_208_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_209_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_210_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_211_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_212_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_213_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_214_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_215_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_216_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_217_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_218_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_219_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_220_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_221_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_222_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_223_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_224_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_225_ ;
 wire net501;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_227_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_228_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_229_ ;
 wire net500;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_231_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_232_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_233_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_234_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_235_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_236_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_237_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_238_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_239_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_240_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_241_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_242_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_243_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_244_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_245_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_246_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_247_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_248_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_249_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_250_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_251_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_252_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_253_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_254_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_255_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_256_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_257_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_258_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_259_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_260_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_261_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_262_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_263_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_264_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_265_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_266_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_267_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_268_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_269_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_270_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_271_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_272_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_273_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_274_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_275_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_276_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_277_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_278_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_279_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_280_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_281_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_282_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_283_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_284_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_285_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_286_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_287_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_288_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_289_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_290_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_291_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_292_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_293_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_294_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_295_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_296_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_297_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_298_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_299_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_300_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_301_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_302_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_303_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_304_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_305_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_306_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_307_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_308_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_309_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_310_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_311_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_312_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_313_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_314_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_315_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_316_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_317_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_318_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_319_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_320_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_321_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_322_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_323_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_324_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_325_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_326_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_327_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_328_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_329_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_330_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_331_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_332_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_333_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_334_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_335_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_336_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_337_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_338_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_339_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_340_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_341_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_342_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_343_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_344_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_345_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_346_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_347_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_348_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_349_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_350_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_351_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_352_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_353_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_354_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_355_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_356_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_357_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_358_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_359_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_360_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_361_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_362_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_363_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_364_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_365_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_366_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_367_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_368_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_369_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_370_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_371_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_372_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_373_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_374_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_375_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_376_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_377_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_378_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_379_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_380_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_381_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_382_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_383_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_384_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_385_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_386_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_387_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_388_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_389_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_390_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_391_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_392_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_393_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_394_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_395_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_396_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_397_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_398_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_399_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_400_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_401_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_402_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_403_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_404_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_405_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_406_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_407_ ;
 wire net546;
 wire net545;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_410_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_411_ ;
 wire net544;
 wire net543;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_414_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_415_ ;
 wire net542;
 wire net541;
 wire net540;
 wire net539;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_420_ ;
 wire net538;
 wire net537;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_423_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_424_ ;
 wire net536;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_426_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_427_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_428_ ;
 wire net535;
 wire net534;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_431_ ;
 wire net533;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_433_ ;
 wire net532;
 wire net531;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_436_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_437_ ;
 wire \i_ibex/if_stage_i/compressed_decoder_i/_438_ ;
 wire net530;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_000_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_001_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_002_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_003_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_004_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_005_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_006_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_007_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_008_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_009_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_010_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_011_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_012_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_013_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_014_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_015_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_016_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_017_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_018_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_019_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_020_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_021_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_022_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_023_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_024_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_025_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_026_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_027_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_028_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_029_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_030_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_031_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_032_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_033_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_034_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_035_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_036_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_037_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_038_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_039_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_040_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_041_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_042_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_043_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_044_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_045_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_046_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_047_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_048_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_049_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_050_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_051_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_052_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_053_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_054_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_055_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_056_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_057_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_058_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_059_ ;
 wire net499;
 wire net498;
 wire net497;
 wire net496;
 wire net495;
 wire net494;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_066_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_067_ ;
 wire net493;
 wire net492;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_070_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_071_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_072_ ;
 wire net491;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_074_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_075_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_076_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_077_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_078_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_079_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_080_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_081_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_082_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_083_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_084_ ;
 wire net490;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_086_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_087_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_088_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_089_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_090_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_091_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_092_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_093_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_094_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_095_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_096_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_097_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_098_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_099_ ;
 wire net489;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_101_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_102_ ;
 wire net488;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_104_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_105_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_106_ ;
 wire net487;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_108_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_109_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_110_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_111_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_112_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_113_ ;
 wire net486;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_115_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_116_ ;
 wire net485;
 wire net484;
 wire net483;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_120_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_121_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_122_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_123_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_124_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_125_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_126_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_127_ ;
 wire net482;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_129_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_130_ ;
 wire net481;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_132_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_133_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_134_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_135_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_136_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_137_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_138_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_139_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_140_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_141_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_142_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_143_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_144_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_145_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_146_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_147_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_148_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_149_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_150_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_151_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_152_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_153_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_154_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_155_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_156_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_157_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_158_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_159_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_160_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_161_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_162_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_163_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_164_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_165_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_166_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_167_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_168_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_169_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_170_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_171_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_172_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_173_ ;
 wire net480;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_175_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_176_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_177_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_178_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_179_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_180_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_181_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_182_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_183_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_184_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_185_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_186_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_187_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_188_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_189_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_190_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_191_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_192_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_193_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_194_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_195_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_196_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_197_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_198_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_199_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_200_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_201_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_202_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_203_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_204_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_205_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_206_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_207_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_208_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_209_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_210_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_211_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_212_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_213_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_214_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_215_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_216_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_217_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_218_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_219_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_220_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_221_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_222_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_223_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_224_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_225_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_226_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_227_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_228_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_229_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_230_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_231_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_232_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_233_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_234_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_235_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_236_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_237_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_238_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_239_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_240_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_241_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_242_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_243_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_244_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_245_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_246_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_247_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_248_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_249_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_250_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_251_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_252_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_253_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_254_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_255_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_256_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_257_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_258_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_259_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_260_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_261_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_262_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_263_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_264_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_265_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_266_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_267_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_268_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_269_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_270_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_271_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_272_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_273_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_274_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_275_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_276_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_277_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_278_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_279_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_280_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_281_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_282_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_283_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_284_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_285_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_286_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_287_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_288_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_289_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_290_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_291_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_292_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_293_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_294_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_295_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_296_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_297_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_298_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_299_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_300_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_301_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_302_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_303_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_304_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_305_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_306_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_307_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_308_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_309_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_310_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_311_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_312_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_313_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_314_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_315_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_316_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_317_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_318_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_319_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_320_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_321_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_322_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_323_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_324_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_325_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_326_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_327_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_328_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_329_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_330_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_331_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_332_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_333_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_334_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_335_ ;
 wire net479;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_337_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_338_ ;
 wire net478;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_340_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_341_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_342_ ;
 wire net477;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_344_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_345_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_346_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_347_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_348_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_349_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_350_ ;
 wire net476;
 wire net475;
 wire net474;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_354_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_355_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_356_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_357_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_358_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_359_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_360_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_361_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_362_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_363_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_364_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_365_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_366_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_367_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_368_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_369_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_370_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_371_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_372_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_373_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_374_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_375_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_376_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_377_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_378_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_379_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_380_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_381_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_382_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_383_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_384_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_385_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_386_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_387_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_388_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_389_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_390_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_391_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_392_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_393_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_394_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_395_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_396_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_397_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_398_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_399_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_400_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_401_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_402_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_403_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_404_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_405_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_406_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_407_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_408_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_409_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_410_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_411_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_412_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_413_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_414_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_415_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/_416_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/discard_req_d ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/discard_req_q ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid_$_AND__Y_B ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__A_B ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__Y_B ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/valid_req_d ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/valid_req_q ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_000_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_001_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_002_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_003_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_004_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_005_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_006_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_007_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_008_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_009_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_010_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_011_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_012_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_013_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_014_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_015_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_016_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_017_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_018_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_019_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_020_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_021_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_022_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_023_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_024_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_025_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_026_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_027_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_028_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_029_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_030_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_031_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_032_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_033_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_034_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_035_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_036_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_037_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_038_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_039_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_040_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_041_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_042_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_043_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_044_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_045_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_046_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_047_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_048_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_049_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_050_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_051_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_052_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_053_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_054_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_055_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_056_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_057_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_058_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_059_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_060_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_061_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_062_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_063_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_064_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_065_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_066_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_067_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_068_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_069_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_070_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_071_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_072_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_073_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_074_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_075_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_076_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_077_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_078_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_079_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_080_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_081_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_082_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_083_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_084_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_085_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_086_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_087_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_088_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_089_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_090_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_091_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_092_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_093_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_094_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_095_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_096_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_097_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_098_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_099_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_100_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_101_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_102_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_103_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_104_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_105_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_106_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_107_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_108_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_109_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_110_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_111_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_112_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_113_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_114_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_115_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_116_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_117_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_118_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_119_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_120_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_121_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_122_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_123_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_124_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_125_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_126_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_127_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_128_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_129_ ;
 wire net473;
 wire net472;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_132_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_133_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_134_ ;
 wire net471;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_136_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_137_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_138_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_139_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_140_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_141_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_142_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_143_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_144_ ;
 wire net470;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_146_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_147_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_149_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_150_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_151_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_152_ ;
 wire net469;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_154_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_155_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ;
 wire net468;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_158_ ;
 wire net467;
 wire net466;
 wire net465;
 wire net464;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_163_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_164_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_165_ ;
 wire net463;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_167_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_168_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_169_ ;
 wire net462;
 wire net461;
 wire net460;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_173_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_174_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_175_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_176_ ;
 wire net459;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_178_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_179_ ;
 wire net458;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_181_ ;
 wire net457;
 wire net456;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_184_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_185_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_186_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_187_ ;
 wire net455;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_189_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_190_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_192_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_193_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_194_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_195_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_196_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_197_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_198_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_199_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_200_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_201_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_202_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_203_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_204_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_205_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_206_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_207_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_208_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_209_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_210_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_211_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_212_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_213_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_214_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_215_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_217_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_218_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_219_ ;
 wire net454;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_221_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_222_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_223_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_224_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ;
 wire net453;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_227_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_228_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_229_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_230_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_231_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_232_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_233_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_234_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_235_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_236_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_237_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_238_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_239_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_240_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_241_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_242_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_243_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_244_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_245_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_246_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_247_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_248_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_249_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_250_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_251_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_252_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_253_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_254_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_255_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_256_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_257_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_258_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_259_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_260_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_261_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_262_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_263_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_264_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_265_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_266_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_267_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_268_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_269_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_270_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_271_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_272_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_273_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_274_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_275_ ;
 wire net452;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_277_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_278_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_279_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_280_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_281_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_282_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_283_ ;
 wire net451;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_285_ ;
 wire net450;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_287_ ;
 wire net449;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_289_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_290_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_291_ ;
 wire net448;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_293_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_294_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_295_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_296_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_297_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_298_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_299_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_300_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_301_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_302_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_303_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_304_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_305_ ;
 wire net447;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_307_ ;
 wire net446;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_309_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_310_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_311_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_312_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_313_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_314_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_315_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_316_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_317_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_318_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_319_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_320_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_321_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_322_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_323_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_324_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_325_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_326_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_327_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_328_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_329_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_330_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_331_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_332_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_333_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_334_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_335_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_336_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_337_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_338_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_339_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_340_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_341_ ;
 wire net445;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_343_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_344_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_345_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_346_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_347_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_348_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_349_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_350_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_351_ ;
 wire net444;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_353_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_354_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_355_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_356_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_357_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_358_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_359_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_360_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_361_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_362_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_363_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_364_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_365_ ;
 wire net443;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_367_ ;
 wire net442;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_369_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_370_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_371_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_372_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_373_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_374_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_375_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_376_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_377_ ;
 wire net441;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_379_ ;
 wire net440;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_381_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_382_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_383_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_384_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_385_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_386_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_387_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_388_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_389_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_390_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_391_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_392_ ;
 wire net439;
 wire net438;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_395_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_396_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_397_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_398_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_399_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_400_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_401_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_402_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_403_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_404_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_405_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_406_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_407_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_408_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_409_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_410_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_411_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_412_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_413_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_414_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_415_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_416_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_417_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_418_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_419_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_420_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_421_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_422_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_423_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_424_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_425_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_426_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_427_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_428_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_429_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_430_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_431_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_432_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_433_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_434_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_435_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_436_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_437_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_438_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_439_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_440_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_441_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_442_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_443_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_444_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_445_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_446_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_447_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_448_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_449_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_450_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_451_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_452_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_453_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_454_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_455_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_456_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_457_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_458_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_459_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_460_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_461_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_462_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_463_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_464_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_465_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_466_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_467_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_468_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_469_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_470_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_471_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_472_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_473_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_474_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_475_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_476_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_477_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_478_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_479_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_480_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_481_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_482_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_483_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_484_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_485_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_486_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_487_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_488_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_489_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_490_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_491_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_492_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_493_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_494_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_495_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_496_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_497_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_498_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_499_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_500_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_501_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_502_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_503_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_504_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_505_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_506_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_507_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_508_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_509_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_510_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_511_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_512_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_513_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_514_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_515_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_516_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_517_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_518_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_519_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_520_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_521_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_522_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_523_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_524_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_525_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_526_ ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_plus2_$_AND__Y_B ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry_$_AND__Y_1_A ;
 wire \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry_$_AND__Y_A ;
 wire \i_ibex/load_store_unit_i/_0000_ ;
 wire \i_ibex/load_store_unit_i/_0001_ ;
 wire \i_ibex/load_store_unit_i/_0002_ ;
 wire \i_ibex/load_store_unit_i/_0003_ ;
 wire \i_ibex/load_store_unit_i/_0004_ ;
 wire \i_ibex/load_store_unit_i/_0005_ ;
 wire \i_ibex/load_store_unit_i/_0006_ ;
 wire \i_ibex/load_store_unit_i/_0007_ ;
 wire \i_ibex/load_store_unit_i/_0008_ ;
 wire \i_ibex/load_store_unit_i/_0009_ ;
 wire \i_ibex/load_store_unit_i/_0010_ ;
 wire \i_ibex/load_store_unit_i/_0011_ ;
 wire \i_ibex/load_store_unit_i/_0012_ ;
 wire \i_ibex/load_store_unit_i/_0013_ ;
 wire \i_ibex/load_store_unit_i/_0014_ ;
 wire \i_ibex/load_store_unit_i/_0015_ ;
 wire \i_ibex/load_store_unit_i/_0016_ ;
 wire \i_ibex/load_store_unit_i/_0017_ ;
 wire \i_ibex/load_store_unit_i/_0018_ ;
 wire \i_ibex/load_store_unit_i/_0019_ ;
 wire \i_ibex/load_store_unit_i/_0020_ ;
 wire \i_ibex/load_store_unit_i/_0021_ ;
 wire \i_ibex/load_store_unit_i/_0022_ ;
 wire \i_ibex/load_store_unit_i/_0023_ ;
 wire \i_ibex/load_store_unit_i/_0024_ ;
 wire \i_ibex/load_store_unit_i/_0025_ ;
 wire \i_ibex/load_store_unit_i/_0026_ ;
 wire \i_ibex/load_store_unit_i/_0027_ ;
 wire \i_ibex/load_store_unit_i/_0028_ ;
 wire \i_ibex/load_store_unit_i/_0029_ ;
 wire \i_ibex/load_store_unit_i/_0030_ ;
 wire \i_ibex/load_store_unit_i/_0031_ ;
 wire \i_ibex/load_store_unit_i/_0032_ ;
 wire \i_ibex/load_store_unit_i/_0033_ ;
 wire \i_ibex/load_store_unit_i/_0034_ ;
 wire \i_ibex/load_store_unit_i/_0035_ ;
 wire \i_ibex/load_store_unit_i/_0036_ ;
 wire \i_ibex/load_store_unit_i/_0037_ ;
 wire \i_ibex/load_store_unit_i/_0038_ ;
 wire \i_ibex/load_store_unit_i/_0039_ ;
 wire \i_ibex/load_store_unit_i/_0040_ ;
 wire \i_ibex/load_store_unit_i/_0041_ ;
 wire \i_ibex/load_store_unit_i/_0042_ ;
 wire \i_ibex/load_store_unit_i/_0043_ ;
 wire \i_ibex/load_store_unit_i/_0044_ ;
 wire \i_ibex/load_store_unit_i/_0045_ ;
 wire \i_ibex/load_store_unit_i/_0046_ ;
 wire \i_ibex/load_store_unit_i/_0047_ ;
 wire \i_ibex/load_store_unit_i/_0048_ ;
 wire \i_ibex/load_store_unit_i/_0049_ ;
 wire \i_ibex/load_store_unit_i/_0050_ ;
 wire \i_ibex/load_store_unit_i/_0051_ ;
 wire \i_ibex/load_store_unit_i/_0052_ ;
 wire \i_ibex/load_store_unit_i/_0053_ ;
 wire \i_ibex/load_store_unit_i/_0054_ ;
 wire \i_ibex/load_store_unit_i/_0055_ ;
 wire \i_ibex/load_store_unit_i/_0056_ ;
 wire \i_ibex/load_store_unit_i/_0057_ ;
 wire \i_ibex/load_store_unit_i/_0058_ ;
 wire \i_ibex/load_store_unit_i/_0059_ ;
 wire \i_ibex/load_store_unit_i/_0060_ ;
 wire \i_ibex/load_store_unit_i/_0061_ ;
 wire \i_ibex/load_store_unit_i/_0062_ ;
 wire \i_ibex/load_store_unit_i/_0063_ ;
 wire \i_ibex/load_store_unit_i/_0064_ ;
 wire \i_ibex/load_store_unit_i/_0065_ ;
 wire \i_ibex/load_store_unit_i/_0066_ ;
 wire \i_ibex/load_store_unit_i/_0067_ ;
 wire net437;
 wire \i_ibex/load_store_unit_i/_0069_ ;
 wire net436;
 wire net435;
 wire \i_ibex/load_store_unit_i/_0072_ ;
 wire \i_ibex/load_store_unit_i/_0073_ ;
 wire net434;
 wire \i_ibex/load_store_unit_i/_0075_ ;
 wire net433;
 wire net432;
 wire \i_ibex/load_store_unit_i/_0078_ ;
 wire net431;
 wire \i_ibex/load_store_unit_i/_0080_ ;
 wire net430;
 wire \i_ibex/load_store_unit_i/_0082_ ;
 wire \i_ibex/load_store_unit_i/_0083_ ;
 wire \i_ibex/load_store_unit_i/_0084_ ;
 wire \i_ibex/load_store_unit_i/_0085_ ;
 wire \i_ibex/load_store_unit_i/_0086_ ;
 wire \i_ibex/load_store_unit_i/_0087_ ;
 wire \i_ibex/load_store_unit_i/_0088_ ;
 wire \i_ibex/load_store_unit_i/_0089_ ;
 wire \i_ibex/load_store_unit_i/_0090_ ;
 wire \i_ibex/load_store_unit_i/_0091_ ;
 wire \i_ibex/load_store_unit_i/_0092_ ;
 wire \i_ibex/load_store_unit_i/_0093_ ;
 wire \i_ibex/load_store_unit_i/_0094_ ;
 wire \i_ibex/load_store_unit_i/_0095_ ;
 wire \i_ibex/load_store_unit_i/_0096_ ;
 wire \i_ibex/load_store_unit_i/_0097_ ;
 wire \i_ibex/load_store_unit_i/_0098_ ;
 wire net429;
 wire net428;
 wire net427;
 wire net426;
 wire \i_ibex/load_store_unit_i/_0103_ ;
 wire net425;
 wire \i_ibex/load_store_unit_i/_0105_ ;
 wire net424;
 wire \i_ibex/load_store_unit_i/_0107_ ;
 wire \i_ibex/load_store_unit_i/_0108_ ;
 wire \i_ibex/load_store_unit_i/_0109_ ;
 wire \i_ibex/load_store_unit_i/_0110_ ;
 wire \i_ibex/load_store_unit_i/_0111_ ;
 wire \i_ibex/load_store_unit_i/_0112_ ;
 wire \i_ibex/load_store_unit_i/_0113_ ;
 wire \i_ibex/load_store_unit_i/_0114_ ;
 wire \i_ibex/load_store_unit_i/_0115_ ;
 wire \i_ibex/load_store_unit_i/_0116_ ;
 wire \i_ibex/load_store_unit_i/_0117_ ;
 wire \i_ibex/load_store_unit_i/_0118_ ;
 wire \i_ibex/load_store_unit_i/_0119_ ;
 wire \i_ibex/load_store_unit_i/_0120_ ;
 wire \i_ibex/load_store_unit_i/_0121_ ;
 wire \i_ibex/load_store_unit_i/_0122_ ;
 wire \i_ibex/load_store_unit_i/_0123_ ;
 wire \i_ibex/load_store_unit_i/_0124_ ;
 wire \i_ibex/load_store_unit_i/_0125_ ;
 wire \i_ibex/load_store_unit_i/_0126_ ;
 wire \i_ibex/load_store_unit_i/_0127_ ;
 wire \i_ibex/load_store_unit_i/_0128_ ;
 wire \i_ibex/load_store_unit_i/_0129_ ;
 wire \i_ibex/load_store_unit_i/_0130_ ;
 wire \i_ibex/load_store_unit_i/_0131_ ;
 wire net423;
 wire net422;
 wire \i_ibex/load_store_unit_i/_0134_ ;
 wire \i_ibex/load_store_unit_i/_0135_ ;
 wire \i_ibex/load_store_unit_i/_0136_ ;
 wire \i_ibex/load_store_unit_i/_0137_ ;
 wire \i_ibex/load_store_unit_i/_0138_ ;
 wire \i_ibex/load_store_unit_i/_0139_ ;
 wire \i_ibex/load_store_unit_i/_0140_ ;
 wire \i_ibex/load_store_unit_i/_0141_ ;
 wire \i_ibex/load_store_unit_i/_0142_ ;
 wire \i_ibex/load_store_unit_i/_0143_ ;
 wire net421;
 wire \i_ibex/load_store_unit_i/_0145_ ;
 wire \i_ibex/load_store_unit_i/_0146_ ;
 wire \i_ibex/load_store_unit_i/_0147_ ;
 wire \i_ibex/load_store_unit_i/_0148_ ;
 wire \i_ibex/load_store_unit_i/_0149_ ;
 wire \i_ibex/load_store_unit_i/_0150_ ;
 wire \i_ibex/load_store_unit_i/_0151_ ;
 wire \i_ibex/load_store_unit_i/_0152_ ;
 wire net420;
 wire \i_ibex/load_store_unit_i/_0154_ ;
 wire \i_ibex/load_store_unit_i/_0155_ ;
 wire net419;
 wire \i_ibex/load_store_unit_i/_0157_ ;
 wire \i_ibex/load_store_unit_i/_0158_ ;
 wire \i_ibex/load_store_unit_i/_0159_ ;
 wire \i_ibex/load_store_unit_i/_0160_ ;
 wire \i_ibex/load_store_unit_i/_0161_ ;
 wire net418;
 wire \i_ibex/load_store_unit_i/_0163_ ;
 wire \i_ibex/load_store_unit_i/_0164_ ;
 wire \i_ibex/load_store_unit_i/_0165_ ;
 wire \i_ibex/load_store_unit_i/_0166_ ;
 wire \i_ibex/load_store_unit_i/_0167_ ;
 wire \i_ibex/load_store_unit_i/_0168_ ;
 wire \i_ibex/load_store_unit_i/_0169_ ;
 wire \i_ibex/load_store_unit_i/_0170_ ;
 wire \i_ibex/load_store_unit_i/_0171_ ;
 wire \i_ibex/load_store_unit_i/_0172_ ;
 wire \i_ibex/load_store_unit_i/_0173_ ;
 wire \i_ibex/load_store_unit_i/_0174_ ;
 wire \i_ibex/load_store_unit_i/_0175_ ;
 wire \i_ibex/load_store_unit_i/_0176_ ;
 wire \i_ibex/load_store_unit_i/_0177_ ;
 wire \i_ibex/load_store_unit_i/_0178_ ;
 wire \i_ibex/load_store_unit_i/_0179_ ;
 wire \i_ibex/load_store_unit_i/_0180_ ;
 wire \i_ibex/load_store_unit_i/_0181_ ;
 wire \i_ibex/load_store_unit_i/_0182_ ;
 wire \i_ibex/load_store_unit_i/_0183_ ;
 wire \i_ibex/load_store_unit_i/_0184_ ;
 wire \i_ibex/load_store_unit_i/_0185_ ;
 wire \i_ibex/load_store_unit_i/_0186_ ;
 wire \i_ibex/load_store_unit_i/_0187_ ;
 wire \i_ibex/load_store_unit_i/_0188_ ;
 wire \i_ibex/load_store_unit_i/_0189_ ;
 wire \i_ibex/load_store_unit_i/_0190_ ;
 wire \i_ibex/load_store_unit_i/_0191_ ;
 wire \i_ibex/load_store_unit_i/_0192_ ;
 wire \i_ibex/load_store_unit_i/_0193_ ;
 wire \i_ibex/load_store_unit_i/_0194_ ;
 wire \i_ibex/load_store_unit_i/_0195_ ;
 wire \i_ibex/load_store_unit_i/_0196_ ;
 wire \i_ibex/load_store_unit_i/_0197_ ;
 wire \i_ibex/load_store_unit_i/_0198_ ;
 wire \i_ibex/load_store_unit_i/_0199_ ;
 wire \i_ibex/load_store_unit_i/_0200_ ;
 wire \i_ibex/load_store_unit_i/_0201_ ;
 wire \i_ibex/load_store_unit_i/_0202_ ;
 wire \i_ibex/load_store_unit_i/_0203_ ;
 wire \i_ibex/load_store_unit_i/_0204_ ;
 wire \i_ibex/load_store_unit_i/_0205_ ;
 wire \i_ibex/load_store_unit_i/_0206_ ;
 wire \i_ibex/load_store_unit_i/_0207_ ;
 wire \i_ibex/load_store_unit_i/_0208_ ;
 wire net417;
 wire net416;
 wire \i_ibex/load_store_unit_i/_0211_ ;
 wire net415;
 wire net414;
 wire net413;
 wire \i_ibex/load_store_unit_i/_0215_ ;
 wire \i_ibex/load_store_unit_i/_0216_ ;
 wire net412;
 wire net411;
 wire \i_ibex/load_store_unit_i/_0219_ ;
 wire net410;
 wire net409;
 wire \i_ibex/load_store_unit_i/_0222_ ;
 wire net408;
 wire net407;
 wire \i_ibex/load_store_unit_i/_0225_ ;
 wire \i_ibex/load_store_unit_i/_0226_ ;
 wire \i_ibex/load_store_unit_i/_0227_ ;
 wire \i_ibex/load_store_unit_i/_0228_ ;
 wire \i_ibex/load_store_unit_i/_0229_ ;
 wire \i_ibex/load_store_unit_i/_0230_ ;
 wire \i_ibex/load_store_unit_i/_0231_ ;
 wire \i_ibex/load_store_unit_i/_0232_ ;
 wire \i_ibex/load_store_unit_i/_0233_ ;
 wire \i_ibex/load_store_unit_i/_0234_ ;
 wire \i_ibex/load_store_unit_i/_0235_ ;
 wire \i_ibex/load_store_unit_i/_0236_ ;
 wire net406;
 wire \i_ibex/load_store_unit_i/_0238_ ;
 wire \i_ibex/load_store_unit_i/_0239_ ;
 wire \i_ibex/load_store_unit_i/_0240_ ;
 wire \i_ibex/load_store_unit_i/_0241_ ;
 wire \i_ibex/load_store_unit_i/_0242_ ;
 wire \i_ibex/load_store_unit_i/_0243_ ;
 wire \i_ibex/load_store_unit_i/_0244_ ;
 wire net405;
 wire net404;
 wire net403;
 wire net402;
 wire \i_ibex/load_store_unit_i/_0249_ ;
 wire \i_ibex/load_store_unit_i/_0250_ ;
 wire \i_ibex/load_store_unit_i/_0251_ ;
 wire net401;
 wire \i_ibex/load_store_unit_i/_0253_ ;
 wire \i_ibex/load_store_unit_i/_0254_ ;
 wire \i_ibex/load_store_unit_i/_0255_ ;
 wire \i_ibex/load_store_unit_i/_0256_ ;
 wire \i_ibex/load_store_unit_i/_0257_ ;
 wire \i_ibex/load_store_unit_i/_0258_ ;
 wire \i_ibex/load_store_unit_i/_0259_ ;
 wire \i_ibex/load_store_unit_i/_0260_ ;
 wire \i_ibex/load_store_unit_i/_0261_ ;
 wire \i_ibex/load_store_unit_i/_0262_ ;
 wire \i_ibex/load_store_unit_i/_0263_ ;
 wire \i_ibex/load_store_unit_i/_0264_ ;
 wire \i_ibex/load_store_unit_i/_0265_ ;
 wire \i_ibex/load_store_unit_i/_0266_ ;
 wire \i_ibex/load_store_unit_i/_0267_ ;
 wire \i_ibex/load_store_unit_i/_0268_ ;
 wire \i_ibex/load_store_unit_i/_0269_ ;
 wire \i_ibex/load_store_unit_i/_0270_ ;
 wire net400;
 wire \i_ibex/load_store_unit_i/_0272_ ;
 wire \i_ibex/load_store_unit_i/_0273_ ;
 wire \i_ibex/load_store_unit_i/_0274_ ;
 wire \i_ibex/load_store_unit_i/_0275_ ;
 wire net399;
 wire net398;
 wire \i_ibex/load_store_unit_i/_0278_ ;
 wire net397;
 wire \i_ibex/load_store_unit_i/_0280_ ;
 wire net396;
 wire \i_ibex/load_store_unit_i/_0282_ ;
 wire \i_ibex/load_store_unit_i/_0283_ ;
 wire \i_ibex/load_store_unit_i/_0284_ ;
 wire \i_ibex/load_store_unit_i/_0285_ ;
 wire \i_ibex/load_store_unit_i/_0286_ ;
 wire \i_ibex/load_store_unit_i/_0287_ ;
 wire \i_ibex/load_store_unit_i/_0288_ ;
 wire \i_ibex/load_store_unit_i/_0289_ ;
 wire \i_ibex/load_store_unit_i/_0290_ ;
 wire \i_ibex/load_store_unit_i/_0291_ ;
 wire \i_ibex/load_store_unit_i/_0292_ ;
 wire \i_ibex/load_store_unit_i/_0293_ ;
 wire \i_ibex/load_store_unit_i/_0294_ ;
 wire \i_ibex/load_store_unit_i/_0295_ ;
 wire \i_ibex/load_store_unit_i/_0296_ ;
 wire \i_ibex/load_store_unit_i/_0297_ ;
 wire \i_ibex/load_store_unit_i/_0298_ ;
 wire \i_ibex/load_store_unit_i/_0299_ ;
 wire \i_ibex/load_store_unit_i/_0300_ ;
 wire \i_ibex/load_store_unit_i/_0301_ ;
 wire \i_ibex/load_store_unit_i/_0302_ ;
 wire net395;
 wire \i_ibex/load_store_unit_i/_0304_ ;
 wire \i_ibex/load_store_unit_i/_0305_ ;
 wire \i_ibex/load_store_unit_i/_0306_ ;
 wire \i_ibex/load_store_unit_i/_0307_ ;
 wire \i_ibex/load_store_unit_i/_0308_ ;
 wire \i_ibex/load_store_unit_i/_0309_ ;
 wire \i_ibex/load_store_unit_i/_0310_ ;
 wire \i_ibex/load_store_unit_i/_0311_ ;
 wire \i_ibex/load_store_unit_i/_0312_ ;
 wire \i_ibex/load_store_unit_i/_0313_ ;
 wire \i_ibex/load_store_unit_i/_0314_ ;
 wire \i_ibex/load_store_unit_i/_0315_ ;
 wire \i_ibex/load_store_unit_i/_0316_ ;
 wire \i_ibex/load_store_unit_i/_0317_ ;
 wire \i_ibex/load_store_unit_i/_0318_ ;
 wire \i_ibex/load_store_unit_i/_0319_ ;
 wire \i_ibex/load_store_unit_i/_0320_ ;
 wire \i_ibex/load_store_unit_i/_0321_ ;
 wire \i_ibex/load_store_unit_i/_0322_ ;
 wire \i_ibex/load_store_unit_i/_0323_ ;
 wire \i_ibex/load_store_unit_i/_0324_ ;
 wire \i_ibex/load_store_unit_i/_0325_ ;
 wire \i_ibex/load_store_unit_i/_0326_ ;
 wire net394;
 wire \i_ibex/load_store_unit_i/_0328_ ;
 wire \i_ibex/load_store_unit_i/_0329_ ;
 wire \i_ibex/load_store_unit_i/_0330_ ;
 wire \i_ibex/load_store_unit_i/_0331_ ;
 wire \i_ibex/load_store_unit_i/_0332_ ;
 wire \i_ibex/load_store_unit_i/_0333_ ;
 wire \i_ibex/load_store_unit_i/_0334_ ;
 wire \i_ibex/load_store_unit_i/_0335_ ;
 wire \i_ibex/load_store_unit_i/_0336_ ;
 wire \i_ibex/load_store_unit_i/_0337_ ;
 wire \i_ibex/load_store_unit_i/_0338_ ;
 wire \i_ibex/load_store_unit_i/_0339_ ;
 wire \i_ibex/load_store_unit_i/_0340_ ;
 wire net393;
 wire \i_ibex/load_store_unit_i/_0342_ ;
 wire \i_ibex/load_store_unit_i/_0343_ ;
 wire \i_ibex/load_store_unit_i/_0344_ ;
 wire \i_ibex/load_store_unit_i/_0345_ ;
 wire \i_ibex/load_store_unit_i/_0346_ ;
 wire \i_ibex/load_store_unit_i/_0347_ ;
 wire net392;
 wire net391;
 wire \i_ibex/load_store_unit_i/_0350_ ;
 wire \i_ibex/load_store_unit_i/_0351_ ;
 wire \i_ibex/load_store_unit_i/_0352_ ;
 wire \i_ibex/load_store_unit_i/_0353_ ;
 wire \i_ibex/load_store_unit_i/_0354_ ;
 wire \i_ibex/load_store_unit_i/_0355_ ;
 wire \i_ibex/load_store_unit_i/_0356_ ;
 wire \i_ibex/load_store_unit_i/_0357_ ;
 wire \i_ibex/load_store_unit_i/_0358_ ;
 wire \i_ibex/load_store_unit_i/_0359_ ;
 wire \i_ibex/load_store_unit_i/_0360_ ;
 wire \i_ibex/load_store_unit_i/_0361_ ;
 wire \i_ibex/load_store_unit_i/_0362_ ;
 wire \i_ibex/load_store_unit_i/_0363_ ;
 wire \i_ibex/load_store_unit_i/_0364_ ;
 wire \i_ibex/load_store_unit_i/_0365_ ;
 wire \i_ibex/load_store_unit_i/_0366_ ;
 wire \i_ibex/load_store_unit_i/_0367_ ;
 wire \i_ibex/load_store_unit_i/_0368_ ;
 wire \i_ibex/load_store_unit_i/_0369_ ;
 wire \i_ibex/load_store_unit_i/_0370_ ;
 wire \i_ibex/load_store_unit_i/_0371_ ;
 wire \i_ibex/load_store_unit_i/_0372_ ;
 wire \i_ibex/load_store_unit_i/_0373_ ;
 wire \i_ibex/load_store_unit_i/_0374_ ;
 wire \i_ibex/load_store_unit_i/_0375_ ;
 wire \i_ibex/load_store_unit_i/_0376_ ;
 wire \i_ibex/load_store_unit_i/_0377_ ;
 wire \i_ibex/load_store_unit_i/_0378_ ;
 wire \i_ibex/load_store_unit_i/_0379_ ;
 wire \i_ibex/load_store_unit_i/_0380_ ;
 wire \i_ibex/load_store_unit_i/_0381_ ;
 wire \i_ibex/load_store_unit_i/_0382_ ;
 wire \i_ibex/load_store_unit_i/_0383_ ;
 wire \i_ibex/load_store_unit_i/_0384_ ;
 wire \i_ibex/load_store_unit_i/_0385_ ;
 wire \i_ibex/load_store_unit_i/_0386_ ;
 wire \i_ibex/load_store_unit_i/_0387_ ;
 wire \i_ibex/load_store_unit_i/_0388_ ;
 wire \i_ibex/load_store_unit_i/_0389_ ;
 wire \i_ibex/load_store_unit_i/_0390_ ;
 wire \i_ibex/load_store_unit_i/_0391_ ;
 wire \i_ibex/load_store_unit_i/_0392_ ;
 wire \i_ibex/load_store_unit_i/_0393_ ;
 wire \i_ibex/load_store_unit_i/_0394_ ;
 wire \i_ibex/load_store_unit_i/_0395_ ;
 wire \i_ibex/load_store_unit_i/_0396_ ;
 wire \i_ibex/load_store_unit_i/_0397_ ;
 wire \i_ibex/load_store_unit_i/_0398_ ;
 wire \i_ibex/load_store_unit_i/_0399_ ;
 wire \i_ibex/load_store_unit_i/_0400_ ;
 wire \i_ibex/load_store_unit_i/_0401_ ;
 wire \i_ibex/load_store_unit_i/_0402_ ;
 wire \i_ibex/load_store_unit_i/_0403_ ;
 wire \i_ibex/load_store_unit_i/_0404_ ;
 wire \i_ibex/load_store_unit_i/_0405_ ;
 wire \i_ibex/load_store_unit_i/_0406_ ;
 wire \i_ibex/load_store_unit_i/_0407_ ;
 wire \i_ibex/load_store_unit_i/_0408_ ;
 wire \i_ibex/load_store_unit_i/_0409_ ;
 wire \i_ibex/load_store_unit_i/_0410_ ;
 wire \i_ibex/load_store_unit_i/_0411_ ;
 wire \i_ibex/load_store_unit_i/_0412_ ;
 wire \i_ibex/load_store_unit_i/_0413_ ;
 wire \i_ibex/load_store_unit_i/_0414_ ;
 wire \i_ibex/load_store_unit_i/_0415_ ;
 wire \i_ibex/load_store_unit_i/_0416_ ;
 wire \i_ibex/load_store_unit_i/_0417_ ;
 wire \i_ibex/load_store_unit_i/_0418_ ;
 wire \i_ibex/load_store_unit_i/_0419_ ;
 wire \i_ibex/load_store_unit_i/_0420_ ;
 wire \i_ibex/load_store_unit_i/_0421_ ;
 wire \i_ibex/load_store_unit_i/_0422_ ;
 wire \i_ibex/load_store_unit_i/_0423_ ;
 wire \i_ibex/load_store_unit_i/_0424_ ;
 wire \i_ibex/load_store_unit_i/_0425_ ;
 wire \i_ibex/load_store_unit_i/_0426_ ;
 wire \i_ibex/load_store_unit_i/_0427_ ;
 wire \i_ibex/load_store_unit_i/_0428_ ;
 wire \i_ibex/load_store_unit_i/_0429_ ;
 wire \i_ibex/load_store_unit_i/_0430_ ;
 wire net390;
 wire net389;
 wire \i_ibex/load_store_unit_i/_0433_ ;
 wire \i_ibex/load_store_unit_i/_0434_ ;
 wire \i_ibex/load_store_unit_i/_0435_ ;
 wire \i_ibex/load_store_unit_i/_0436_ ;
 wire \i_ibex/load_store_unit_i/_0437_ ;
 wire \i_ibex/load_store_unit_i/_0438_ ;
 wire \i_ibex/load_store_unit_i/_0439_ ;
 wire \i_ibex/load_store_unit_i/_0440_ ;
 wire \i_ibex/load_store_unit_i/_0441_ ;
 wire \i_ibex/load_store_unit_i/_0442_ ;
 wire \i_ibex/load_store_unit_i/_0443_ ;
 wire \i_ibex/load_store_unit_i/_0444_ ;
 wire \i_ibex/load_store_unit_i/_0445_ ;
 wire \i_ibex/load_store_unit_i/_0446_ ;
 wire \i_ibex/load_store_unit_i/_0447_ ;
 wire \i_ibex/load_store_unit_i/_0448_ ;
 wire \i_ibex/load_store_unit_i/_0449_ ;
 wire \i_ibex/load_store_unit_i/_0450_ ;
 wire \i_ibex/load_store_unit_i/_0451_ ;
 wire \i_ibex/load_store_unit_i/_0452_ ;
 wire \i_ibex/load_store_unit_i/_0453_ ;
 wire \i_ibex/load_store_unit_i/_0454_ ;
 wire \i_ibex/load_store_unit_i/_0455_ ;
 wire \i_ibex/load_store_unit_i/_0456_ ;
 wire \i_ibex/load_store_unit_i/_0457_ ;
 wire \i_ibex/load_store_unit_i/_0458_ ;
 wire \i_ibex/load_store_unit_i/_0459_ ;
 wire \i_ibex/load_store_unit_i/_0460_ ;
 wire \i_ibex/load_store_unit_i/_0461_ ;
 wire \i_ibex/load_store_unit_i/_0462_ ;
 wire \i_ibex/load_store_unit_i/_0463_ ;
 wire \i_ibex/load_store_unit_i/_0464_ ;
 wire \i_ibex/load_store_unit_i/_0465_ ;
 wire \i_ibex/load_store_unit_i/_0466_ ;
 wire \i_ibex/load_store_unit_i/_0467_ ;
 wire \i_ibex/load_store_unit_i/_0468_ ;
 wire \i_ibex/load_store_unit_i/_0469_ ;
 wire \i_ibex/load_store_unit_i/_0470_ ;
 wire \i_ibex/load_store_unit_i/_0471_ ;
 wire \i_ibex/load_store_unit_i/_0472_ ;
 wire \i_ibex/load_store_unit_i/_0473_ ;
 wire \i_ibex/load_store_unit_i/_0474_ ;
 wire \i_ibex/load_store_unit_i/_0475_ ;
 wire \i_ibex/load_store_unit_i/_0476_ ;
 wire \i_ibex/load_store_unit_i/_0477_ ;
 wire \i_ibex/load_store_unit_i/_0478_ ;
 wire \i_ibex/load_store_unit_i/_0479_ ;
 wire \i_ibex/load_store_unit_i/_0480_ ;
 wire \i_ibex/load_store_unit_i/_0481_ ;
 wire \i_ibex/load_store_unit_i/_0482_ ;
 wire \i_ibex/load_store_unit_i/_0483_ ;
 wire \i_ibex/load_store_unit_i/_0484_ ;
 wire \i_ibex/load_store_unit_i/_0485_ ;
 wire \i_ibex/load_store_unit_i/_0486_ ;
 wire \i_ibex/load_store_unit_i/_0487_ ;
 wire \i_ibex/load_store_unit_i/_0488_ ;
 wire \i_ibex/load_store_unit_i/_0489_ ;
 wire \i_ibex/load_store_unit_i/_0490_ ;
 wire \i_ibex/load_store_unit_i/_0491_ ;
 wire \i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ;
 wire \i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ;
 wire \i_ibex/load_store_unit_i/data_sign_ext_q ;
 wire \i_ibex/load_store_unit_i/data_type_q_$_NOT__A_1_Y ;
 wire \i_ibex/load_store_unit_i/data_type_q_$_NOT__A_Y ;
 wire \i_ibex/load_store_unit_i/data_we_q ;
 wire \i_ibex/load_store_unit_i/handle_misaligned_q ;
 wire \i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg_E_$_AND__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ;
 wire \i_ibex/load_store_unit_i/lsu_err_q ;
 wire \i_ibex/load_store_unit_i/lsu_err_q_$_NOT__A_Y ;
 wire \i_ibex/load_store_unit_i/lsu_rdata_valid_o_$_AND__Y_B ;
 wire \i_ibex/load_store_unit_i/pmp_err_q ;
 wire \i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_1_Y ;
 wire \i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ;
 wire \i_ibex/wb_i/_000_ ;
 wire net388;
 wire net387;
 wire net386;
 wire \i_ibex/wb_i/_004_ ;
 wire \i_ibex/wb_i/_005_ ;
 wire \i_ibex/wb_i/_006_ ;
 wire \i_ibex/wb_i/_007_ ;
 wire \i_ibex/wb_i/_008_ ;
 wire \i_ibex/wb_i/_009_ ;
 wire \i_ibex/wb_i/_010_ ;
 wire \i_ibex/wb_i/_011_ ;
 wire \i_ibex/wb_i/_012_ ;
 wire net385;
 wire \i_ibex/wb_i/_014_ ;
 wire net384;
 wire \i_ibex/wb_i/_016_ ;
 wire \i_ibex/wb_i/_017_ ;
 wire \i_ibex/wb_i/_018_ ;
 wire \i_ibex/wb_i/_019_ ;
 wire \i_ibex/wb_i/_020_ ;
 wire \i_ibex/wb_i/_021_ ;
 wire \i_ibex/wb_i/_022_ ;
 wire \i_ibex/wb_i/_023_ ;
 wire \i_ibex/wb_i/_024_ ;
 wire net383;
 wire \i_ibex/wb_i/_026_ ;
 wire net382;
 wire \i_ibex/wb_i/_028_ ;
 wire \i_ibex/wb_i/_029_ ;
 wire \i_ibex/wb_i/_030_ ;
 wire \i_ibex/wb_i/_031_ ;
 wire \i_ibex/wb_i/_032_ ;
 wire \i_ibex/wb_i/_033_ ;
 wire \i_ibex/wb_i/_034_ ;
 wire \i_ibex/wb_i/_035_ ;
 wire \i_ibex/wb_i/_036_ ;
 wire \i_ibex/wb_i/_037_ ;
 wire \i_ibex/wb_i/_038_ ;
 wire \i_ibex/wb_i/_039_ ;
 wire VDD;
 wire VSS;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net43;
 wire net44;
 wire net45;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire clk_i_regs;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_leaf_0_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_24_clk_i_regs;
 wire clknet_leaf_25_clk_i_regs;
 wire clknet_leaf_27_clk_i_regs;
 wire clknet_leaf_28_clk_i_regs;
 wire clknet_leaf_29_clk_i_regs;
 wire clknet_leaf_30_clk_i_regs;
 wire clknet_leaf_31_clk_i_regs;
 wire clknet_leaf_32_clk_i_regs;
 wire clknet_leaf_33_clk_i_regs;
 wire clknet_leaf_34_clk_i_regs;
 wire clknet_leaf_35_clk_i_regs;
 wire clknet_leaf_36_clk_i_regs;
 wire clknet_leaf_37_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire clknet_leaf_39_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire clknet_leaf_41_clk_i_regs;
 wire clknet_leaf_42_clk_i_regs;
 wire clknet_leaf_43_clk_i_regs;
 wire clknet_leaf_45_clk_i_regs;
 wire clknet_leaf_46_clk_i_regs;
 wire clknet_leaf_47_clk_i_regs;
 wire clknet_leaf_48_clk_i_regs;
 wire clknet_leaf_49_clk_i_regs;
 wire clknet_leaf_50_clk_i_regs;
 wire clknet_leaf_51_clk_i_regs;
 wire clknet_leaf_52_clk_i_regs;
 wire clknet_leaf_53_clk_i_regs;
 wire clknet_leaf_54_clk_i_regs;
 wire clknet_leaf_55_clk_i_regs;
 wire clknet_leaf_56_clk_i_regs;
 wire clknet_leaf_57_clk_i_regs;
 wire clknet_leaf_58_clk_i_regs;
 wire clknet_leaf_59_clk_i_regs;
 wire clknet_leaf_60_clk_i_regs;
 wire clknet_leaf_61_clk_i_regs;
 wire clknet_leaf_62_clk_i_regs;
 wire clknet_leaf_63_clk_i_regs;
 wire clknet_leaf_64_clk_i_regs;
 wire clknet_leaf_65_clk_i_regs;
 wire clknet_leaf_66_clk_i_regs;
 wire clknet_leaf_67_clk_i_regs;
 wire clknet_leaf_68_clk_i_regs;
 wire clknet_leaf_69_clk_i_regs;
 wire clknet_leaf_70_clk_i_regs;
 wire clknet_leaf_71_clk_i_regs;
 wire clknet_leaf_72_clk_i_regs;
 wire clknet_leaf_73_clk_i_regs;
 wire clknet_leaf_74_clk_i_regs;
 wire clknet_leaf_75_clk_i_regs;
 wire clknet_leaf_76_clk_i_regs;
 wire clknet_leaf_77_clk_i_regs;
 wire clknet_leaf_78_clk_i_regs;
 wire clknet_leaf_79_clk_i_regs;
 wire clknet_leaf_80_clk_i_regs;
 wire clknet_leaf_81_clk_i_regs;
 wire clknet_leaf_82_clk_i_regs;
 wire clknet_leaf_83_clk_i_regs;
 wire clknet_leaf_84_clk_i_regs;
 wire clknet_leaf_85_clk_i_regs;
 wire clknet_leaf_86_clk_i_regs;
 wire clknet_leaf_87_clk_i_regs;
 wire clknet_leaf_88_clk_i_regs;
 wire clknet_leaf_89_clk_i_regs;
 wire clknet_leaf_91_clk_i_regs;
 wire clknet_leaf_92_clk_i_regs;
 wire clknet_leaf_93_clk_i_regs;
 wire clknet_leaf_94_clk_i_regs;
 wire clknet_leaf_95_clk_i_regs;
 wire clknet_leaf_96_clk_i_regs;
 wire clknet_leaf_97_clk_i_regs;
 wire clknet_leaf_98_clk_i_regs;
 wire clknet_leaf_99_clk_i_regs;
 wire clknet_leaf_103_clk_i_regs;
 wire clknet_leaf_104_clk_i_regs;
 wire clknet_leaf_105_clk_i_regs;
 wire clknet_leaf_106_clk_i_regs;
 wire clknet_leaf_107_clk_i_regs;
 wire clknet_leaf_108_clk_i_regs;
 wire clknet_leaf_109_clk_i_regs;
 wire clknet_leaf_110_clk_i_regs;
 wire clknet_leaf_111_clk_i_regs;
 wire clknet_leaf_112_clk_i_regs;
 wire clknet_leaf_113_clk_i_regs;
 wire clknet_leaf_114_clk_i_regs;
 wire clknet_leaf_115_clk_i_regs;
 wire clknet_leaf_116_clk_i_regs;
 wire clknet_leaf_117_clk_i_regs;
 wire clknet_leaf_118_clk_i_regs;
 wire clknet_leaf_119_clk_i_regs;
 wire clknet_leaf_120_clk_i_regs;
 wire clknet_leaf_121_clk_i_regs;
 wire clknet_leaf_122_clk_i_regs;
 wire clknet_leaf_123_clk_i_regs;
 wire clknet_leaf_124_clk_i_regs;
 wire clknet_leaf_125_clk_i_regs;
 wire clknet_leaf_126_clk_i_regs;
 wire clknet_leaf_128_clk_i_regs;
 wire clknet_leaf_129_clk_i_regs;
 wire clknet_leaf_130_clk_i_regs;
 wire clknet_leaf_131_clk_i_regs;
 wire clknet_leaf_132_clk_i_regs;
 wire clknet_leaf_133_clk_i_regs;
 wire clknet_leaf_134_clk_i_regs;
 wire clknet_leaf_135_clk_i_regs;
 wire clknet_leaf_137_clk_i_regs;
 wire clknet_leaf_138_clk_i_regs;
 wire clknet_leaf_139_clk_i_regs;
 wire clknet_leaf_140_clk_i_regs;
 wire clknet_leaf_141_clk_i_regs;
 wire clknet_leaf_142_clk_i_regs;
 wire clknet_leaf_143_clk_i_regs;
 wire clknet_leaf_144_clk_i_regs;
 wire clknet_leaf_145_clk_i_regs;
 wire clknet_leaf_146_clk_i_regs;
 wire clknet_leaf_147_clk_i_regs;
 wire clknet_leaf_148_clk_i_regs;
 wire clknet_leaf_149_clk_i_regs;
 wire clknet_leaf_150_clk_i_regs;
 wire clknet_leaf_151_clk_i_regs;
 wire clknet_leaf_152_clk_i_regs;
 wire clknet_leaf_153_clk_i_regs;
 wire clknet_leaf_154_clk_i_regs;
 wire clknet_leaf_155_clk_i_regs;
 wire clknet_leaf_156_clk_i_regs;
 wire clknet_leaf_157_clk_i_regs;
 wire clknet_leaf_158_clk_i_regs;
 wire clknet_leaf_159_clk_i_regs;
 wire clknet_leaf_160_clk_i_regs;
 wire clknet_leaf_161_clk_i_regs;
 wire clknet_leaf_162_clk_i_regs;
 wire clknet_leaf_163_clk_i_regs;
 wire clknet_0_clk_i_regs;
 wire clknet_4_0_0_clk_i_regs;
 wire clknet_4_1_0_clk_i_regs;
 wire clknet_4_2_0_clk_i_regs;
 wire clknet_4_3_0_clk_i_regs;
 wire clknet_4_4_0_clk_i_regs;
 wire clknet_4_5_0_clk_i_regs;
 wire clknet_4_6_0_clk_i_regs;
 wire clknet_4_7_0_clk_i_regs;
 wire clknet_4_8_0_clk_i_regs;
 wire clknet_4_9_0_clk_i_regs;
 wire clknet_4_10_0_clk_i_regs;
 wire clknet_4_11_0_clk_i_regs;
 wire clknet_4_12_0_clk_i_regs;
 wire clknet_4_13_0_clk_i_regs;
 wire clknet_4_14_0_clk_i_regs;
 wire clknet_4_15_0_clk_i_regs;
 wire clknet_5_0__leaf_clk_i_regs;
 wire clknet_5_1__leaf_clk_i_regs;
 wire clknet_5_2__leaf_clk_i_regs;
 wire clknet_5_3__leaf_clk_i_regs;
 wire clknet_5_4__leaf_clk_i_regs;
 wire clknet_5_5__leaf_clk_i_regs;
 wire clknet_5_6__leaf_clk_i_regs;
 wire clknet_5_7__leaf_clk_i_regs;
 wire clknet_5_8__leaf_clk_i_regs;
 wire clknet_5_9__leaf_clk_i_regs;
 wire clknet_5_10__leaf_clk_i_regs;
 wire clknet_5_11__leaf_clk_i_regs;
 wire clknet_5_12__leaf_clk_i_regs;
 wire clknet_5_13__leaf_clk_i_regs;
 wire clknet_5_14__leaf_clk_i_regs;
 wire clknet_5_15__leaf_clk_i_regs;
 wire clknet_5_16__leaf_clk_i_regs;
 wire clknet_5_17__leaf_clk_i_regs;
 wire clknet_5_18__leaf_clk_i_regs;
 wire clknet_5_19__leaf_clk_i_regs;
 wire clknet_5_20__leaf_clk_i_regs;
 wire clknet_5_21__leaf_clk_i_regs;
 wire clknet_5_22__leaf_clk_i_regs;
 wire clknet_5_23__leaf_clk_i_regs;
 wire clknet_5_24__leaf_clk_i_regs;
 wire clknet_5_25__leaf_clk_i_regs;
 wire clknet_5_26__leaf_clk_i_regs;
 wire clknet_5_27__leaf_clk_i_regs;
 wire clknet_5_28__leaf_clk_i_regs;
 wire clknet_5_29__leaf_clk_i_regs;
 wire clknet_5_30__leaf_clk_i_regs;
 wire clknet_5_31__leaf_clk_i_regs;
 wire delaynet_0_clk_sys;
 wire delaynet_1_clk_sys;
 wire delaynet_2_clk_sys;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire [31:0] \i_ibex/alu_adder_result_ex ;
 wire [31:0] \i_ibex/alu_operand_a_ex ;
 wire [31:0] \i_ibex/alu_operand_b_ex ;
 wire [6:0] \i_ibex/alu_operator_ex ;
 wire [31:0] \i_ibex/branch_target_ex ;
 wire [31:0] \i_ibex/cs_registers_i/csr_wdata_int ;
 wire [31:0] \i_ibex/cs_registers_i/dcsr_d ;
 wire [31:0] \i_ibex/cs_registers_i/dcsr_q ;
 wire [31:0] \i_ibex/cs_registers_i/depc_d ;
 wire [31:0] \i_ibex/cs_registers_i/dscratch0_q ;
 wire [31:0] \i_ibex/cs_registers_i/dscratch1_q ;
 wire [31:0] \i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value ;
 wire [194:0] \i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y ;
 wire [6:0] \i_ibex/cs_registers_i/mcause_d ;
 wire [6:0] \i_ibex/cs_registers_i/mcause_q ;
 wire [0:0] \i_ibex/cs_registers_i/mcycle_counter_i/counter_upd ;
 wire [31:0] \i_ibex/cs_registers_i/mepc_d ;
 wire [2047:0] \i_ibex/cs_registers_i/mhpmcounter ;
 wire [2:0] \i_ibex/cs_registers_i/mhpmcounter_we ;
 wire [2:0] \i_ibex/cs_registers_i/mhpmcounterh_we ;
 wire [18:0] \i_ibex/cs_registers_i/mie_q ;
 wire [63:0] \i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o ;
 wire [63:0] \i_ibex/cs_registers_i/minstret_raw ;
 wire [31:0] \i_ibex/cs_registers_i/mscratch_q ;
 wire [6:0] \i_ibex/cs_registers_i/mstack_cause_q ;
 wire [31:0] \i_ibex/cs_registers_i/mstack_epc_q ;
 wire [2:0] \i_ibex/cs_registers_i/mstack_q ;
 wire [5:0] \i_ibex/cs_registers_i/mstatus_d ;
 wire [4:0] \i_ibex/cs_registers_i/mstatus_q ;
 wire [31:0] \i_ibex/cs_registers_i/mtval_d ;
 wire [31:0] \i_ibex/cs_registers_i/mtval_q ;
 wire [31:0] \i_ibex/cs_registers_i/mtvec_d ;
 wire [11:0] \i_ibex/csr_addr ;
 wire [31:0] \i_ibex/csr_depc ;
 wire [31:0] \i_ibex/csr_mepc ;
 wire [31:0] \i_ibex/csr_mtval ;
 wire [31:0] \i_ibex/csr_mtvec ;
 wire [1:0] \i_ibex/csr_op ;
 wire [135:0] \i_ibex/csr_pmp_addr ;
 wire [23:0] \i_ibex/csr_pmp_cfg ;
 wire [1:0] \i_ibex/csr_pmp_mseccfg ;
 wire [31:0] \i_ibex/csr_rdata ;
 wire [2:0] \i_ibex/debug_cause ;
 wire [33:0] \i_ibex/ex_block_i/alu_adder_result_ext ;
 wire [6:0] \i_ibex/exc_cause ;
 wire [1:0] \i_ibex/exc_pc_mux_id ;
 wire [1:0] \i_ibex/g_no_pmp.unused_priv_lvl_ls ;
 wire [1:0] \i_ibex/id_stage_i/alu_op_a_mux_sel_dec ;
 wire [3:0] \i_ibex/id_stage_i/controller_i/ctrl_fsm_cs ;
 wire [2:0] \i_ibex/id_stage_i/imm_b_mux_sel_dec ;
 wire [31:0] \i_ibex/id_stage_i/imm_b_type ;
 wire [31:0] \i_ibex/id_stage_i/imm_i_type ;
 wire [31:0] \i_ibex/id_stage_i/imm_j_type ;
 wire [31:0] \i_ibex/id_stage_i/imm_s_type ;
 wire [31:0] \i_ibex/id_stage_i/imm_u_type ;
 wire [31:0] \i_ibex/id_stage_i/zimm_rs1_type ;
 wire [31:0] \i_ibex/if_stage_i/fetch_addr_n ;
 wire [31:0] \i_ibex/if_stage_i/fetch_rdata ;
 wire [31:0] \i_ibex/if_stage_i/instr_decompressed ;
 wire [1:0] \i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q ;
 wire [1:0] \i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_s ;
 wire [31:0] \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q ;
 wire [1:0] \i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy ;
 wire [2:0] \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q ;
 wire [0:0] \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry ;
 wire [95:0] \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q ;
 wire [2:0] \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d ;
 wire [0:0] \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_q ;
 wire [1:0] \i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q ;
 wire [1:0] \i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_s ;
 wire [31:0] \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q ;
 wire [66:0] \i_ibex/imd_val_d_ex ;
 wire [67:0] \i_ibex/imd_val_q_ex ;
 wire [0:0] \i_ibex/imd_val_we_ex ;
 wire [31:0] \i_ibex/instr_rdata_alu_id ;
 wire [15:0] \i_ibex/instr_rdata_c_id ;
 wire [31:0] \i_ibex/instr_rdata_id ;
 wire [18:0] \i_ibex/irqs ;
 wire [3:0] \i_ibex/load_store_unit_i/data_be_o_$_MUX__Y_A ;
 wire [1:0] \i_ibex/load_store_unit_i/data_type_q ;
 wire [2:0] \i_ibex/load_store_unit_i/ls_fsm_cs ;
 wire [1:0] \i_ibex/load_store_unit_i/rdata_offset_q ;
 wire [23:0] \i_ibex/load_store_unit_i/rdata_q ;
 wire [31:0] \i_ibex/lsu_addr_last ;
 wire [1:0] \i_ibex/lsu_type ;
 wire [31:0] \i_ibex/lsu_wdata ;
 wire [31:0] \i_ibex/multdiv_operand_a_ex ;
 wire [31:0] \i_ibex/multdiv_operand_b_ex ;
 wire [1:0] \i_ibex/multdiv_operator_ex ;
 wire [1:0] \i_ibex/multdiv_signed_mode_ex ;
 wire [31:0] \i_ibex/pc_id ;
 wire [31:0] \i_ibex/pc_if ;
 wire [2:0] \i_ibex/pc_mux_id ;
 wire [1:0] \i_ibex/priv_mode_id ;
 wire [31:0] \i_ibex/result_ex ;
 wire [4:0] \i_ibex/rf_raddr_a ;
 wire [4:0] \i_ibex/rf_raddr_b ;
 wire [31:0] \i_ibex/rf_rdata_a ;
 wire [31:0] \i_ibex/rf_rdata_b ;
 wire [4:0] \i_ibex/rf_waddr_id ;
 wire [4:0] \i_ibex/rf_waddr_wb ;
 wire [31:0] \i_ibex/rf_wdata_id ;
 wire [31:0] \i_ibex/rf_wdata_lsu ;
 wire [31:0] \i_ibex/rf_wdata_wb ;

 sg13g2_tielo \i_ibex/if_stage_i/_735__42  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net42));
 sg13g2_or3_2 \i_ibex/_02_  (.A(\i_ibex/lsu_busy ),
    .B(\i_ibex/ctrl_busy ),
    .C(\i_ibex/if_busy ),
    .X(core_busy_o),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/_03_  (.A(\i_ibex/alu_operand_b_ex [11]),
    .B(net617),
    .X(\i_ibex/csr_addr [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(net1049),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_05_  (.A(net617),
    .B(\i_ibex/alu_operand_b_ex [10]),
    .X(\i_ibex/csr_addr [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_06_  (.A(net617),
    .B(\i_ibex/alu_operand_b_ex [1]),
    .X(\i_ibex/csr_addr [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_07_  (.A(net617),
    .B(net490),
    .X(\i_ibex/csr_addr [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/_08_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [9]),
    .X(\i_ibex/csr_addr [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/_09_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [8]),
    .X(\i_ibex/csr_addr [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_10_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [7]),
    .X(\i_ibex/csr_addr [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_11_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [6]),
    .X(\i_ibex/csr_addr [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/_12_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [5]),
    .X(\i_ibex/csr_addr [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_13_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [4]),
    .X(\i_ibex/csr_addr [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/_14_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [3]),
    .X(\i_ibex/csr_addr [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/_15_  (.A(net616),
    .B(\i_ibex/alu_operand_b_ex [2]),
    .X(\i_ibex/csr_addr [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/_16_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/lsu_resp_err ),
    .B(\i_ibex/lsu_store_err ),
    .A(\i_ibex/lsu_load_err ));
 sg13g2_nor2b_1 \i_ibex/_17_  (.A(net707),
    .B_N(\i_ibex/id_in_ready ),
    .Y(\i_ibex/perf_iside_wait ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_3__46  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net46));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net474),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(net1046),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1044 (.A(net1045),
    .X(net1044),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1134_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0010_ ),
    .B(net1089),
    .A(net1091));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(net1045),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(\i_ibex/cs_registers_i/_0025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/cs_registers_i/_1137_  (.Y(\i_ibex/cs_registers_i/_0013_ ),
    .A(net588),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1041 (.A(net1042),
    .X(net1041),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(\i_ibex/cs_registers_i/_0026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1140_  (.Y(\i_ibex/cs_registers_i/_0016_ ),
    .A(net1068),
    .B(net506),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1141_  (.Y(\i_ibex/cs_registers_i/_0017_ ),
    .A(net1061),
    .B(\i_ibex/cs_registers_i/_0016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1039 (.A(\i_ibex/cs_registers_i/_0054_ ),
    .X(net1039),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1144_  (.B1(\i_ibex/csr_addr [5]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0020_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0010_ ),
    .A2(\i_ibex/cs_registers_i/_0017_ ));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1036 (.A(net1038),
    .X(net1036),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/cs_registers_i/_1147_  (.A(\i_ibex/csr_addr [5]),
    .B(net1067),
    .C(net506),
    .D(\i_ibex/cs_registers_i/_0010_ ),
    .X(\i_ibex/cs_registers_i/_0023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(\i_ibex/cs_registers_i/_0054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1149_  (.A(net586),
    .B(net1089),
    .Y(\i_ibex/cs_registers_i/_0025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1150_  (.A(net1065),
    .B(net518),
    .Y(\i_ibex/cs_registers_i/_0026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1151_  (.Y(\i_ibex/cs_registers_i/_0027_ ),
    .A(net1041),
    .B(net1040),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/cs_registers_i/_1152_  (.A(\i_ibex/csr_addr [5]),
    .B(net1092),
    .C(\i_ibex/cs_registers_i/_0027_ ),
    .X(\i_ibex/cs_registers_i/_0028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1034 (.A(net1035),
    .X(net1034),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(\i_ibex/cs_registers_i/_0078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(net1033),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1156_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0032_ ),
    .A(\i_ibex/csr_addr [7]),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1157_  (.Y(\i_ibex/cs_registers_i/_0033_ ),
    .A(\i_ibex/csr_addr [9]),
    .B(\i_ibex/csr_addr [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1031 (.X(net1031),
    .A(\i_ibex/cs_registers_i/_0086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1030 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_084_ ),
    .X(net1030),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1160_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0036_ ),
    .B(\i_ibex/csr_addr [11]),
    .A(net1106));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1161_  (.A(\i_ibex/cs_registers_i/_0033_ ),
    .B(\i_ibex/cs_registers_i/_0036_ ),
    .Y(\i_ibex/cs_registers_i/_0037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1162_  (.Y(\i_ibex/cs_registers_i/_0038_ ),
    .A(\i_ibex/cs_registers_i/_0032_ ),
    .B(net464),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1163_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1095),
    .C1(\i_ibex/cs_registers_i/_0038_ ),
    .B1(\i_ibex/cs_registers_i/_0028_ ),
    .A1(\i_ibex/cs_registers_i/_0020_ ),
    .Y(\i_ibex/cs_registers_i/_0039_ ),
    .A2(\i_ibex/cs_registers_i/_0023_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1164_  (.A(\i_ibex/csr_addr [9]),
    .B(\i_ibex/csr_addr [8]),
    .X(\i_ibex/cs_registers_i/_0040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1165_  (.A(net1106),
    .B(\i_ibex/csr_addr [11]),
    .Y(\i_ibex/cs_registers_i/_0041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1166_  (.Y(\i_ibex/cs_registers_i/_0042_ ),
    .A(\i_ibex/cs_registers_i/_0040_ ),
    .B(\i_ibex/cs_registers_i/_0041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_1167_  (.Y(\i_ibex/cs_registers_i/_0043_ ),
    .A(net484),
    .B(net1065),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1168_  (.A(net1093),
    .B(net518),
    .C(\i_ibex/cs_registers_i/_0043_ ),
    .Y(\i_ibex/cs_registers_i/_0044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1029 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_102_ ),
    .X(net1029),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1170_  (.A(net1097),
    .B(net1090),
    .C(net588),
    .D(net1088),
    .Y(\i_ibex/cs_registers_i/_0046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/cs_registers_i/_1171_  (.Y(\i_ibex/cs_registers_i/_0047_ ),
    .B(net1062),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net506));
 sg13g2_or4_2 \i_ibex/cs_registers_i/_1172_  (.A(net484),
    .B(net1093),
    .C(net1097),
    .D(net1090),
    .X(\i_ibex/cs_registers_i/_0048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_1173_  (.A(net1061),
    .B(net1088),
    .C(\i_ibex/cs_registers_i/_0047_ ),
    .Y(\i_ibex/cs_registers_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0048_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1174_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0044_ ),
    .A2(net462),
    .Y(\i_ibex/cs_registers_i/_0050_ ),
    .B1(\i_ibex/cs_registers_i/_0049_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1175_  (.A(\i_ibex/cs_registers_i/_0042_ ),
    .B(\i_ibex/cs_registers_i/_0050_ ),
    .Y(\i_ibex/cs_registers_i/_0051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1176_  (.A(net518),
    .B_N(net1068),
    .Y(\i_ibex/cs_registers_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/_1177_  (.B(net588),
    .A(net497),
    .X(\i_ibex/cs_registers_i/_0053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/cs_registers_i/_1178_  (.Y(\i_ibex/cs_registers_i/_0054_ ),
    .A(net1069),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1179_  (.Y(\i_ibex/cs_registers_i/_0055_ ),
    .B1(\i_ibex/cs_registers_i/_0053_ ),
    .B2(net1035),
    .A2(\i_ibex/cs_registers_i/_0052_ ),
    .A1(net1061),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1180_  (.B(\i_ibex/csr_addr [8]),
    .C(net1106),
    .A(\i_ibex/csr_addr [9]),
    .Y(\i_ibex/cs_registers_i/_0056_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net1091));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1181_  (.A(\i_ibex/csr_addr [3]),
    .B(\i_ibex/cs_registers_i/_0056_ ),
    .Y(\i_ibex/cs_registers_i/_0057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1182_  (.Y(\i_ibex/cs_registers_i/_0058_ ),
    .B(\i_ibex/csr_addr [11]),
    .A_N(net483),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1183_  (.A(net1095),
    .B(net1098),
    .C(\i_ibex/cs_registers_i/_0058_ ),
    .Y(\i_ibex/cs_registers_i/_0059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/_1184_  (.B(\i_ibex/cs_registers_i/_0057_ ),
    .C(\i_ibex/cs_registers_i/_0059_ ),
    .Y(\i_ibex/cs_registers_i/_0060_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/cs_registers_i/_0055_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1185_  (.B(\i_ibex/csr_addr [8]),
    .C(net1106),
    .A(\i_ibex/csr_addr [9]),
    .Y(\i_ibex/cs_registers_i/_0061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/_1186_  (.B(net484),
    .C(net1098),
    .Y(\i_ibex/cs_registers_i/_0062_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/csr_addr [11]));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1187_  (.A(net1094),
    .B(net1092),
    .C(\i_ibex/cs_registers_i/_0061_ ),
    .D(\i_ibex/cs_registers_i/_0062_ ),
    .Y(\i_ibex/cs_registers_i/_0063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1188_  (.B(\i_ibex/cs_registers_i/_0016_ ),
    .C(\i_ibex/cs_registers_i/_0063_ ),
    .A(net1041),
    .Y(\i_ibex/cs_registers_i/_0064_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1189_  (.Y(\i_ibex/cs_registers_i/_0065_ ),
    .A(net1061),
    .B(\i_ibex/cs_registers_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1190_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0066_ ),
    .B(net1094),
    .A(net483));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1191_  (.Y(\i_ibex/cs_registers_i/_0067_ ),
    .B(\i_ibex/csr_addr [11]),
    .A_N(net1106),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_1192_  (.A(\i_ibex/cs_registers_i/_0033_ ),
    .B(\i_ibex/cs_registers_i/_0066_ ),
    .C(\i_ibex/cs_registers_i/_0067_ ),
    .Y(\i_ibex/cs_registers_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1193_  (.B1(\i_ibex/cs_registers_i/_0068_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0069_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0010_ ),
    .A2(\i_ibex/cs_registers_i/_0065_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1194_  (.A(net484),
    .B_N(net1093),
    .Y(\i_ibex/cs_registers_i/_0070_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1195_  (.A(net1097),
    .B(net1091),
    .Y(\i_ibex/cs_registers_i/_0071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1196_  (.B(\i_ibex/cs_registers_i/_0041_ ),
    .C(net473),
    .A(\i_ibex/cs_registers_i/_0040_ ),
    .Y(\i_ibex/cs_registers_i/_0072_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0071_ ));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1197_  (.A(net518),
    .B_N(net586),
    .Y(\i_ibex/cs_registers_i/_0073_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1198_  (.A(net588),
    .B_N(net506),
    .Y(\i_ibex/cs_registers_i/_0074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1199_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1035),
    .A2(\i_ibex/cs_registers_i/_0073_ ),
    .Y(\i_ibex/cs_registers_i/_0075_ ),
    .B1(\i_ibex/cs_registers_i/_0074_ ));
 sg13g2_or3_1 \i_ibex/cs_registers_i/_1200_  (.A(\i_ibex/csr_addr [3]),
    .B(\i_ibex/cs_registers_i/_0072_ ),
    .C(\i_ibex/cs_registers_i/_0075_ ),
    .X(\i_ibex/cs_registers_i/_0076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1201_  (.B(\i_ibex/cs_registers_i/_0064_ ),
    .C(\i_ibex/cs_registers_i/_0069_ ),
    .A(\i_ibex/cs_registers_i/_0060_ ),
    .Y(\i_ibex/cs_registers_i/_0077_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0076_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1202_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0078_ ),
    .B(net1088),
    .A(net588));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_1203_  (.A(net1095),
    .B(net1032),
    .C(\i_ibex/cs_registers_i/_0056_ ),
    .Y(\i_ibex/cs_registers_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0062_ ));
 sg13g2_buf_2 fanout1028 (.A(net1029),
    .X(net1028),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1205_  (.Y(\i_ibex/cs_registers_i/_0081_ ),
    .A(net1041),
    .B(\i_ibex/cs_registers_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1206_  (.A(\i_ibex/cs_registers_i/_0081_ ),
    .B(\i_ibex/cs_registers_i/_0072_ ),
    .Y(\i_ibex/cs_registers_i/_0082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1207_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0083_ ),
    .B(\i_ibex/cs_registers_i/_0082_ ),
    .A(net460));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1208_  (.A(\i_ibex/cs_registers_i/_0039_ ),
    .B(\i_ibex/cs_registers_i/_0051_ ),
    .C(\i_ibex/cs_registers_i/_0077_ ),
    .D(\i_ibex/cs_registers_i/_0083_ ),
    .Y(\i_ibex/cs_registers_i/_0084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1027 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_350_ ),
    .X(net1027),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_1210_  (.A(net1065),
    .B(net506),
    .C(net1088),
    .Y(\i_ibex/cs_registers_i/_0086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1211_  (.A(net586),
    .B(net1031),
    .X(\i_ibex/cs_registers_i/_0087_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1026 (.A(net1027),
    .X(net1026),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1025 (.X(net1025),
    .A(net1027),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1024 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_350_ ),
    .X(net1024),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_350_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(\i_ibex/cs_registers_i/_0948_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1021 (.A(\i_ibex/cs_registers_i/_0948_ ),
    .X(net1021),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1218_  (.Y(\i_ibex/cs_registers_i/_0094_ ),
    .A(\i_ibex/csr_mepc [31]),
    .B(net1071),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(net1021),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1019 (.A(net1020),
    .X(net1019),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1221_  (.A0(\i_ibex/cs_registers_i/mcause_q [6]),
    .A1(\i_ibex/cs_registers_i/mtval_q [31]),
    .S(net1067),
    .X(\i_ibex/cs_registers_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1222_  (.Y(\i_ibex/cs_registers_i/_0098_ ),
    .A(net519),
    .B(\i_ibex/cs_registers_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1223_  (.B1(\i_ibex/cs_registers_i/_0098_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0099_ ),
    .VSS(VSS),
    .A1(net507),
    .A2(\i_ibex/cs_registers_i/_0094_ ));
 sg13g2_buf_2 fanout1018 (.A(\i_ibex/ex_block_i/alu_i/_0094_ ),
    .X(net1018),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1225_  (.Y(\i_ibex/cs_registers_i/_0101_ ),
    .B1(\i_ibex/cs_registers_i/_0099_ ),
    .B2(\i_ibex/cs_registers_i/_0025_ ),
    .A2(net456),
    .A1(irqs_i[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1226_  (.Y(\i_ibex/cs_registers_i/_0102_ ),
    .B(net1093),
    .A_N(net483),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1227_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0103_ ),
    .B(net1090),
    .A(net1097));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1228_  (.A(\i_ibex/cs_registers_i/_0033_ ),
    .B(\i_ibex/cs_registers_i/_0036_ ),
    .C(\i_ibex/cs_registers_i/_0102_ ),
    .D(\i_ibex/cs_registers_i/_0103_ ),
    .Y(\i_ibex/cs_registers_i/_0104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1229_  (.Y(\i_ibex/cs_registers_i/_0105_ ),
    .B(net453),
    .A_N(\i_ibex/cs_registers_i/_0101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_1230_  (.A(net1068),
    .B(\i_ibex/cs_registers_i/_0033_ ),
    .C(\i_ibex/cs_registers_i/_0066_ ),
    .Y(\i_ibex/cs_registers_i/_0106_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0067_ ));
 sg13g2_nand2b_2 \i_ibex/cs_registers_i/_1231_  (.Y(\i_ibex/cs_registers_i/_0107_ ),
    .B(net1097),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1090));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1232_  (.A(net1032),
    .B(\i_ibex/cs_registers_i/_0107_ ),
    .Y(\i_ibex/cs_registers_i/_0108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1234_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2047]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [63]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1235_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2015]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [31]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1016 (.A(net1017),
    .X(net1016),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1237_  (.Y(\i_ibex/cs_registers_i/_0113_ ),
    .B1(\i_ibex/cs_registers_i/_0111_ ),
    .B2(net463),
    .A2(\i_ibex/cs_registers_i/_0110_ ),
    .A1(\i_ibex/cs_registers_i/_0108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1238_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0114_ ),
    .A(\i_ibex/cs_registers_i/_0113_ ),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_1239_  (.A(\i_ibex/cs_registers_i/_0033_ ),
    .B(\i_ibex/cs_registers_i/_0036_ ),
    .C(\i_ibex/cs_registers_i/_0048_ ),
    .Y(\i_ibex/cs_registers_i/_0115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1240_  (.A(net457),
    .B(\i_ibex/cs_registers_i/_0115_ ),
    .X(\i_ibex/cs_registers_i/_0116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(net1018),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1242_  (.B(net1040),
    .C(\i_ibex/cs_registers_i/_0071_ ),
    .A(net1041),
    .Y(\i_ibex/cs_registers_i/_0118_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1244_  (.A(net1093),
    .B_N(net484),
    .Y(\i_ibex/cs_registers_i/_0120_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1245_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [31]),
    .A2(\i_ibex/cs_registers_i/_0070_ ),
    .Y(\i_ibex/cs_registers_i/_0121_ ),
    .B1(\i_ibex/cs_registers_i/_0120_ ));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1246_  (.A(\i_ibex/cs_registers_i/_0042_ ),
    .B(\i_ibex/cs_registers_i/_0118_ ),
    .C(\i_ibex/cs_registers_i/_0121_ ),
    .Y(\i_ibex/cs_registers_i/_0122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1247_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/mie_q [15]),
    .C1(\i_ibex/cs_registers_i/_0122_ ),
    .B1(net436),
    .A1(\i_ibex/cs_registers_i/_0106_ ),
    .Y(\i_ibex/cs_registers_i/_0123_ ),
    .A2(\i_ibex/cs_registers_i/_0114_ ));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_1248_  (.A(net1094),
    .B(net1098),
    .C(\i_ibex/cs_registers_i/_0056_ ),
    .Y(\i_ibex/cs_registers_i/_0124_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0058_ ));
 sg13g2_and2_2 \i_ibex/cs_registers_i/_1249_  (.A(net457),
    .B(\i_ibex/cs_registers_i/_0124_ ),
    .X(\i_ibex/cs_registers_i/_0125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_1251_  (.A(net1094),
    .B(\i_ibex/cs_registers_i/_0056_ ),
    .C(\i_ibex/cs_registers_i/_0062_ ),
    .Y(\i_ibex/cs_registers_i/_0127_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1252_  (.A(net1032),
    .B(\i_ibex/cs_registers_i/_0016_ ),
    .Y(\i_ibex/cs_registers_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/cs_registers_i/_1253_  (.A(\i_ibex/cs_registers_i/_0127_ ),
    .B(\i_ibex/cs_registers_i/_0128_ ),
    .X(\i_ibex/cs_registers_i/_0129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(\i_ibex/ex_block_i/alu_i/_0098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1255_  (.Y(\i_ibex/cs_registers_i/_0131_ ),
    .B1(net450),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [31]),
    .A2(net991),
    .A1(net1),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1011 (.A(net1012),
    .X(net1011),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1257_  (.A(net464),
    .B(\i_ibex/cs_registers_i/_0049_ ),
    .X(\i_ibex/cs_registers_i/_0133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1258_  (.Y(\i_ibex/cs_registers_i/_0134_ ),
    .B(net518),
    .A_N(net1066),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1259_  (.A(net1032),
    .B(\i_ibex/cs_registers_i/_0134_ ),
    .Y(\i_ibex/cs_registers_i/_0135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1260_  (.A(\i_ibex/cs_registers_i/_0063_ ),
    .B(\i_ibex/cs_registers_i/_0135_ ),
    .X(\i_ibex/cs_registers_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1010 (.A(\i_ibex/ex_block_i/alu_i/_0098_ ),
    .X(net1010),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1009 (.A(net1010),
    .X(net1009),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1008 (.A(net1009),
    .X(net1008),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1264_  (.A(net1103),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [31]),
    .Y(\i_ibex/cs_registers_i/_0140_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1265_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [31]),
    .A2(net1104),
    .Y(\i_ibex/cs_registers_i/_0141_ ),
    .B1(\i_ibex/cs_registers_i/_0140_ ));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(net1010),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1006 (.A(\i_ibex/cs_registers_i/_0169_ ),
    .X(net1006),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1268_  (.B(net1037),
    .C(net510),
    .A(\i_ibex/cs_registers_i/dscratch0_q [31]),
    .Y(\i_ibex/cs_registers_i/_0144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1269_  (.B1(\i_ibex/cs_registers_i/_0144_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0145_ ),
    .VSS(VSS),
    .A1(net509),
    .A2(\i_ibex/cs_registers_i/_0141_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1270_  (.A(net458),
    .B(\i_ibex/cs_registers_i/_0145_ ),
    .X(\i_ibex/cs_registers_i/_0146_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1271_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [31]),
    .C1(\i_ibex/cs_registers_i/_0146_ ),
    .B1(net446),
    .A1(\i_ibex/csr_mtvec [31]),
    .Y(\i_ibex/cs_registers_i/_0147_ ),
    .A2(net986));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1272_  (.B(\i_ibex/cs_registers_i/_0123_ ),
    .C(\i_ibex/cs_registers_i/_0131_ ),
    .A(\i_ibex/cs_registers_i/_0105_ ),
    .Y(\i_ibex/cs_registers_i/_0148_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0147_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1273_  (.A(net978),
    .B_N(\i_ibex/cs_registers_i/_0148_ ),
    .Y(\i_ibex/csr_rdata [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1274_  (.Y(\i_ibex/cs_registers_i/_0149_ ),
    .A(net690),
    .B(\i_ibex/csr_rdata [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1275_  (.Y(\i_ibex/cs_registers_i/_0150_ ),
    .A(net689),
    .B(\i_ibex/csr_op [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1276_  (.Y(\i_ibex/cs_registers_i/_0151_ ),
    .A(\i_ibex/alu_operand_a_ex [31]),
    .B(net631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1277_  (.B1(\i_ibex/cs_registers_i/_0151_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [31]),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_a_ex [31]),
    .A2(\i_ibex/cs_registers_i/_0149_ ));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(net1006),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/cs_registers_i/_1279_  (.Y(\i_ibex/cs_registers_i/_0153_ ),
    .B(net689),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net979));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(net1005),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(net1006),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1002 (.A(\i_ibex/cs_registers_i/_0188_ ),
    .X(net1002),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1283_  (.S0(net1063),
    .A0(\i_ibex/cs_registers_i/mscratch_q [5]),
    .A1(\i_ibex/csr_mepc [5]),
    .A2(\i_ibex/cs_registers_i/mcause_q [5]),
    .A3(\i_ibex/cs_registers_i/mtval_q [5]),
    .S1(net521),
    .X(\i_ibex/cs_registers_i/_0157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1001 (.A(net1002),
    .X(net1001),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1285_  (.A(net1032),
    .B(\i_ibex/cs_registers_i/_0072_ ),
    .Y(\i_ibex/cs_registers_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_1286_  (.A(net1094),
    .B(\i_ibex/cs_registers_i/_0061_ ),
    .C(\i_ibex/cs_registers_i/_0062_ ),
    .Y(\i_ibex/cs_registers_i/_0160_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/_1287_  (.A(net1090),
    .B(net1041),
    .C(net1040),
    .D(\i_ibex/cs_registers_i/_0160_ ),
    .X(\i_ibex/cs_registers_i/_0161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1289_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0163_ ),
    .A(net1096),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1290_  (.Y(\i_ibex/cs_registers_i/_0164_ ),
    .A(net484),
    .B(\i_ibex/cs_registers_i/_0163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1291_  (.A(\i_ibex/cs_registers_i/_0042_ ),
    .B(\i_ibex/cs_registers_i/_0118_ ),
    .C(\i_ibex/cs_registers_i/_0164_ ),
    .Y(\i_ibex/cs_registers_i/_0165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout999 (.A(\i_ibex/cs_registers_i/_0188_ ),
    .X(net999),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1293_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/dcsr_q [5]),
    .C1(net983),
    .B1(net445),
    .A1(\i_ibex/cs_registers_i/_0157_ ),
    .Y(\i_ibex/cs_registers_i/_0167_ ),
    .A2(\i_ibex/cs_registers_i/_0159_ ));
 sg13g2_buf_2 fanout998 (.A(net999),
    .X(net998),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1295_  (.A(net462),
    .B(\i_ibex/cs_registers_i/_0106_ ),
    .X(\i_ibex/cs_registers_i/_0169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout997 (.A(\i_ibex/ex_block_i/alu_i/_0087_ ),
    .X(net997),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout996 (.A(\i_ibex/ex_block_i/alu_i/_0087_ ),
    .X(net996),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout995 (.A(\i_ibex/ex_block_i/alu_i/_0087_ ),
    .X(net995),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout994 (.A(net995),
    .X(net994),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1300_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1989]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [5]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0174_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1301_  (.Y(\i_ibex/cs_registers_i/_0175_ ),
    .B1(net1003),
    .B2(\i_ibex/cs_registers_i/_0174_ ),
    .A2(net984),
    .A1(\i_ibex/csr_mtvec [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout993 (.A(net994),
    .X(net993),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout992 (.A(net995),
    .X(net992),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout991 (.X(net991),
    .A(\i_ibex/cs_registers_i/_0125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1305_  (.A2(net456),
    .A1(net2),
    .B1(\i_ibex/cs_registers_i/_0135_ ),
    .X(\i_ibex/cs_registers_i/_0179_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1306_  (.Y(\i_ibex/cs_registers_i/_0180_ ),
    .B1(\i_ibex/cs_registers_i/_0124_ ),
    .B2(\i_ibex/cs_registers_i/_0179_ ),
    .A2(net449),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout990 (.A(net991),
    .X(net990),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout989 (.A(\i_ibex/cs_registers_i/_0125_ ),
    .X(net989),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1310_  (.Y(\i_ibex/cs_registers_i/_0184_ ),
    .A(\i_ibex/csr_depc [5]),
    .B(net1063),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1311_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [5]),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [5]),
    .S(net1062),
    .X(\i_ibex/cs_registers_i/_0185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1312_  (.Y(\i_ibex/cs_registers_i/_0186_ ),
    .A(net520),
    .B(\i_ibex/cs_registers_i/_0185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1313_  (.B1(\i_ibex/cs_registers_i/_0186_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0187_ ),
    .VSS(VSS),
    .A1(net511),
    .A2(\i_ibex/cs_registers_i/_0184_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1314_  (.A(\i_ibex/cs_registers_i/_0106_ ),
    .B(\i_ibex/cs_registers_i/_0108_ ),
    .X(\i_ibex/cs_registers_i/_0188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout987 (.A(\i_ibex/cs_registers_i/_0133_ ),
    .X(net987),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout986 (.A(net987),
    .X(net986),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1317_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2021]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [37]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0191_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1318_  (.Y(\i_ibex/cs_registers_i/_0192_ ),
    .B1(net998),
    .B2(\i_ibex/cs_registers_i/_0191_ ),
    .A2(\i_ibex/cs_registers_i/_0187_ ),
    .A1(net459),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1319_  (.A(\i_ibex/cs_registers_i/_0167_ ),
    .B(\i_ibex/cs_registers_i/_0175_ ),
    .C(\i_ibex/cs_registers_i/_0180_ ),
    .D(\i_ibex/cs_registers_i/_0192_ ),
    .X(\i_ibex/cs_registers_i/_0193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1320_  (.A(net547),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0193_ ),
    .Y(\i_ibex/cs_registers_i/_0194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1321_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0194_ ),
    .Y(\i_ibex/cs_registers_i/_0195_ ),
    .A2(net634),
    .A1(net547));
 sg13g2_inv_4 \i_ibex/cs_registers_i/_1322_  (.A(\i_ibex/cs_registers_i/_0195_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1323_  (.Y(\i_ibex/cs_registers_i/_0196_ ),
    .A(\i_ibex/cs_registers_i/_0070_ ),
    .B(\i_ibex/cs_registers_i/_0071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1324_  (.Y(\i_ibex/cs_registers_i/_0197_ ),
    .B(net518),
    .A_N(net586),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout985 (.A(net986),
    .X(net985),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout984 (.A(\i_ibex/cs_registers_i/_0133_ ),
    .X(net984),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1327_  (.A(\i_ibex/cs_registers_i/mtval_q [4]),
    .B(net1063),
    .X(\i_ibex/cs_registers_i/_0200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1328_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcause_q [4]),
    .A2(net1035),
    .Y(\i_ibex/cs_registers_i/_0201_ ),
    .B1(\i_ibex/cs_registers_i/_0200_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1329_  (.A(net1089),
    .B(\i_ibex/cs_registers_i/_0196_ ),
    .C(\i_ibex/cs_registers_i/_0197_ ),
    .D(\i_ibex/cs_registers_i/_0201_ ),
    .Y(\i_ibex/cs_registers_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1330_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [4]),
    .A2(\i_ibex/cs_registers_i/_0070_ ),
    .Y(\i_ibex/cs_registers_i/_0203_ ),
    .B1(\i_ibex/cs_registers_i/_0120_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1331_  (.A(\i_ibex/cs_registers_i/_0118_ ),
    .B(\i_ibex/cs_registers_i/_0203_ ),
    .Y(\i_ibex/cs_registers_i/_0204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout983 (.A(\i_ibex/cs_registers_i/_0165_ ),
    .X(net983),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1333_  (.B1(net466),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0206_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0202_ ),
    .A2(\i_ibex/cs_registers_i/_0204_ ));
 sg13g2_buf_2 fanout982 (.A(net983),
    .X(net982),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1335_  (.Y(\i_ibex/cs_registers_i/_0208_ ),
    .B1(net989),
    .B2(net3),
    .A2(\i_ibex/cs_registers_i/_0082_ ),
    .A1(\i_ibex/csr_mepc [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout981 (.A(\i_ibex/ex_block_i/alu_i/_1021_ ),
    .X(net981),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout980 (.A(\i_ibex/cs_registers_i/_0084_ ),
    .X(net980),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net980),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout978 (.A(net979),
    .X(net978),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1340_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2020]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [36]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0213_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1341_  (.Y(\i_ibex/cs_registers_i/_0214_ ),
    .B1(net998),
    .B2(\i_ibex/cs_registers_i/_0213_ ),
    .A2(net984),
    .A1(\i_ibex/csr_mtvec [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net978),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1343_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [4]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [4]),
    .A2(\i_ibex/csr_depc [4]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [4]),
    .S1(net1100),
    .X(\i_ibex/cs_registers_i/_0216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(net980),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1345_  (.Y(\i_ibex/cs_registers_i/_0218_ ),
    .A(net463),
    .B(\i_ibex/cs_registers_i/_0106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net976),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1347_  (.A(net520),
    .B_N(\i_ibex/cs_registers_i/mhpmcounter [1988]),
    .Y(\i_ibex/cs_registers_i/_0220_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1348_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net521),
    .A2(\i_ibex/cs_registers_i/minstret_raw [4]),
    .Y(\i_ibex/cs_registers_i/_0221_ ),
    .B1(\i_ibex/cs_registers_i/_0220_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1349_  (.A(\i_ibex/cs_registers_i/_0218_ ),
    .B(\i_ibex/cs_registers_i/_0221_ ),
    .Y(\i_ibex/cs_registers_i/_0222_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1350_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net461),
    .C1(\i_ibex/cs_registers_i/_0222_ ),
    .B1(\i_ibex/cs_registers_i/_0216_ ),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [4]),
    .Y(\i_ibex/cs_registers_i/_0223_ ),
    .A2(net447));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1351_  (.B(\i_ibex/cs_registers_i/_0208_ ),
    .C(\i_ibex/cs_registers_i/_0214_ ),
    .A(\i_ibex/cs_registers_i/_0206_ ),
    .Y(\i_ibex/cs_registers_i/_0224_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0223_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1352_  (.A(net975),
    .B_N(\i_ibex/cs_registers_i/_0224_ ),
    .Y(\i_ibex/csr_rdata [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1353_  (.Y(\i_ibex/cs_registers_i/_0225_ ),
    .A(net690),
    .B(\i_ibex/csr_rdata [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout974 (.A(\i_ibex/cs_registers_i/csr_wdata_int [0]),
    .X(net974),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1355_  (.Y(\i_ibex/cs_registers_i/_0227_ ),
    .A(net545),
    .B(net634),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1356_  (.B1(\i_ibex/cs_registers_i/_0227_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [4]),
    .VSS(VSS),
    .A1(net545),
    .A2(\i_ibex/cs_registers_i/_0225_ ));
 sg13g2_and2_2 \i_ibex/cs_registers_i/_1357_  (.A(net689),
    .B(\i_ibex/csr_op [0]),
    .X(\i_ibex/cs_registers_i/_0228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout973 (.X(net973),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout972 (.A(\i_ibex/cs_registers_i/csr_wdata_int [1]),
    .X(net972),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1360_  (.Y(\i_ibex/cs_registers_i/_0231_ ),
    .A(\i_ibex/csr_depc [3]),
    .B(net1067),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1361_  (.B(net1035),
    .C(net507),
    .A(\i_ibex/cs_registers_i/dscratch0_q [3]),
    .Y(\i_ibex/cs_registers_i/_0232_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1362_  (.B1(\i_ibex/cs_registers_i/_0232_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0233_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0231_ ));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1363_  (.A(net507),
    .B(\i_ibex/csr_addr [3]),
    .Y(\i_ibex/cs_registers_i/_0234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout970 (.A(\i_ibex/rf_we_id ),
    .X(net970),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1366_  (.Y(\i_ibex/cs_registers_i/_0237_ ),
    .A(\i_ibex/csr_mepc [3]),
    .B(net1067),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/_1367_  (.B(net589),
    .C(net4),
    .Y(\i_ibex/cs_registers_i/_0238_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1067));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1368_  (.B1(\i_ibex/cs_registers_i/_0238_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0239_ ),
    .VSS(VSS),
    .A1(net590),
    .A2(\i_ibex/cs_registers_i/_0237_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1369_  (.Y(\i_ibex/cs_registers_i/_0240_ ),
    .B1(\i_ibex/cs_registers_i/_0234_ ),
    .B2(\i_ibex/cs_registers_i/_0239_ ),
    .A2(\i_ibex/cs_registers_i/_0128_ ),
    .A1(\i_ibex/cs_registers_i/mtval_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1370_  (.A(\i_ibex/cs_registers_i/_0072_ ),
    .B(\i_ibex/cs_registers_i/_0240_ ),
    .Y(\i_ibex/cs_registers_i/_0241_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1371_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net461),
    .C1(\i_ibex/cs_registers_i/_0241_ ),
    .B1(\i_ibex/cs_registers_i/_0233_ ),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [3]),
    .Y(\i_ibex/cs_registers_i/_0242_ ),
    .A2(net447));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1372_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0243_ ),
    .B(\i_ibex/cs_registers_i/_0107_ ),
    .A(net1032));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1373_  (.A(net520),
    .B_N(\i_ibex/cs_registers_i/mhpmcounter [2019]),
    .Y(\i_ibex/cs_registers_i/_0244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1374_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net519),
    .A2(\i_ibex/cs_registers_i/minstret_raw [35]),
    .Y(\i_ibex/cs_registers_i/_0245_ ),
    .B1(\i_ibex/cs_registers_i/_0244_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1375_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [3]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1376_  (.Y(\i_ibex/cs_registers_i/_0247_ ),
    .A(net463),
    .B(\i_ibex/cs_registers_i/_0246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1377_  (.B1(\i_ibex/cs_registers_i/_0247_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0248_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0243_ ),
    .A2(\i_ibex/cs_registers_i/_0245_ ));
 sg13g2_or3_1 \i_ibex/cs_registers_i/_1378_  (.A(net1106),
    .B(net1097),
    .C(net1065),
    .X(\i_ibex/cs_registers_i/_0249_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1379_  (.B(net1098),
    .C(net1065),
    .A(net1106),
    .Y(\i_ibex/cs_registers_i/_0250_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1380_  (.A(\i_ibex/csr_addr [11]),
    .B_N(net484),
    .Y(\i_ibex/cs_registers_i/_0251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1381_  (.A(net1093),
    .B(net1091),
    .C(net518),
    .Y(\i_ibex/cs_registers_i/_0252_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1382_  (.B(\i_ibex/cs_registers_i/_0040_ ),
    .C(\i_ibex/cs_registers_i/_0251_ ),
    .A(net1041),
    .Y(\i_ibex/cs_registers_i/_0253_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0252_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1383_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0253_ ),
    .Y(\i_ibex/cs_registers_i/_0254_ ),
    .A2(\i_ibex/cs_registers_i/_0250_ ),
    .A1(\i_ibex/cs_registers_i/_0249_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1384_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0106_ ),
    .C1(\i_ibex/cs_registers_i/_0254_ ),
    .B1(\i_ibex/cs_registers_i/_0248_ ),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [3]),
    .Y(\i_ibex/cs_registers_i/_0255_ ),
    .A2(\i_ibex/cs_registers_i/_0129_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1385_  (.Y(\i_ibex/cs_registers_i/_0256_ ),
    .A(net473),
    .B(net462),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1386_  (.A0(\i_ibex/cs_registers_i/mscratch_q [3]),
    .A1(\i_ibex/cs_registers_i/mcause_q [3]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0257_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1387_  (.Y(\i_ibex/cs_registers_i/_0258_ ),
    .A(net1034),
    .B(\i_ibex/cs_registers_i/_0257_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_1388_  (.A(net484),
    .B(net1096),
    .C(net1098),
    .Y(\i_ibex/cs_registers_i/_0259_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net1091));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1389_  (.A0(\i_ibex/csr_mstatus_mie ),
    .A1(\i_ibex/cs_registers_i/mie_q [18]),
    .S(net586),
    .X(\i_ibex/cs_registers_i/_0260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1390_  (.B(net1031),
    .C(\i_ibex/cs_registers_i/_0260_ ),
    .A(\i_ibex/cs_registers_i/_0259_ ),
    .Y(\i_ibex/cs_registers_i/_0261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1391_  (.B1(\i_ibex/cs_registers_i/_0261_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0262_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0256_ ),
    .A2(\i_ibex/cs_registers_i/_0258_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1392_  (.Y(\i_ibex/cs_registers_i/_0263_ ),
    .B1(\i_ibex/cs_registers_i/_0262_ ),
    .B2(net465),
    .A2(net445),
    .A1(\i_ibex/cs_registers_i/dcsr_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1393_  (.Y(\i_ibex/cs_registers_i/_0264_ ),
    .B1(net988),
    .B2(net5),
    .A2(net984),
    .A1(\i_ibex/csr_mtvec [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/_1394_  (.X(\i_ibex/cs_registers_i/_0265_ ),
    .A(\i_ibex/cs_registers_i/_0255_ ),
    .B(\i_ibex/cs_registers_i/_0263_ ),
    .C(\i_ibex/cs_registers_i/_0264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1395_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net975),
    .Y(\i_ibex/csr_rdata [3]),
    .A2(\i_ibex/cs_registers_i/_0265_ ),
    .A1(\i_ibex/cs_registers_i/_0242_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1396_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net689),
    .A2(\i_ibex/csr_rdata [3]),
    .Y(\i_ibex/cs_registers_i/_0266_ ),
    .B1(net543));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1397_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net543),
    .A2(\i_ibex/cs_registers_i/_0228_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [3]),
    .B1(\i_ibex/cs_registers_i/_0266_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1398_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2018]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [34]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0267_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1399_  (.A(net520),
    .B_N(\i_ibex/cs_registers_i/mhpmcounter [1986]),
    .Y(\i_ibex/cs_registers_i/_0268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1400_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net521),
    .A2(\i_ibex/cs_registers_i/minstret_raw [2]),
    .Y(\i_ibex/cs_registers_i/_0269_ ),
    .B1(\i_ibex/cs_registers_i/_0268_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1401_  (.A(\i_ibex/cs_registers_i/_0218_ ),
    .B(\i_ibex/cs_registers_i/_0269_ ),
    .Y(\i_ibex/cs_registers_i/_0270_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1402_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net998),
    .C1(\i_ibex/cs_registers_i/_0270_ ),
    .B1(\i_ibex/cs_registers_i/_0267_ ),
    .A1(\i_ibex/debug_single_step ),
    .Y(\i_ibex/cs_registers_i/_0271_ ),
    .A2(\i_ibex/cs_registers_i/_0161_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1403_  (.A(net473),
    .B(net462),
    .X(\i_ibex/cs_registers_i/_0272_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1404_  (.Y(\i_ibex/cs_registers_i/_0273_ ),
    .A(\i_ibex/csr_mepc [2]),
    .B(net1063),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1405_  (.A0(\i_ibex/cs_registers_i/mcause_q [2]),
    .A1(\i_ibex/cs_registers_i/mtval_q [2]),
    .S(net1063),
    .X(\i_ibex/cs_registers_i/_0274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1406_  (.Y(\i_ibex/cs_registers_i/_0275_ ),
    .A(net519),
    .B(\i_ibex/cs_registers_i/_0274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1407_  (.B1(\i_ibex/cs_registers_i/_0275_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0276_ ),
    .VSS(VSS),
    .A1(net512),
    .A2(\i_ibex/cs_registers_i/_0273_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1408_  (.Y(\i_ibex/cs_registers_i/_0277_ ),
    .B1(\i_ibex/cs_registers_i/_0120_ ),
    .B2(\i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y [194]),
    .A2(net473),
    .A1(\i_ibex/cs_registers_i/mscratch_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1409_  (.A(net1088),
    .B(\i_ibex/cs_registers_i/_0047_ ),
    .C(\i_ibex/cs_registers_i/_0048_ ),
    .Y(\i_ibex/cs_registers_i/_0278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1410_  (.B1(\i_ibex/cs_registers_i/_0278_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0279_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_mtvec [2]),
    .A2(net1061));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1411_  (.B1(\i_ibex/cs_registers_i/_0279_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0280_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0118_ ),
    .A2(\i_ibex/cs_registers_i/_0277_ ));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1412_  (.A2(\i_ibex/cs_registers_i/_0276_ ),
    .A1(\i_ibex/cs_registers_i/_0272_ ),
    .B1(\i_ibex/cs_registers_i/_0280_ ),
    .X(\i_ibex/cs_registers_i/_0281_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1413_  (.Y(\i_ibex/cs_registers_i/_0282_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [2]),
    .B(net509),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/_1414_  (.B(net1068),
    .C(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_control ),
    .Y(\i_ibex/cs_registers_i/_0283_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net512));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1415_  (.B1(\i_ibex/cs_registers_i/_0283_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0284_ ),
    .VSS(VSS),
    .A1(net1068),
    .A2(\i_ibex/cs_registers_i/_0282_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1416_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1041),
    .A2(\i_ibex/cs_registers_i/_0284_ ),
    .Y(\i_ibex/cs_registers_i/_0285_ ),
    .B1(net1090));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1417_  (.A(net1033),
    .B(\i_ibex/cs_registers_i/_0047_ ),
    .Y(\i_ibex/cs_registers_i/_0286_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1418_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0287_ ),
    .A(net1091),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1419_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/dscratch0_q [2]),
    .C1(\i_ibex/cs_registers_i/_0287_ ),
    .B1(\i_ibex/cs_registers_i/_0135_ ),
    .A1(\i_ibex/csr_depc [2]),
    .Y(\i_ibex/cs_registers_i/_0288_ ),
    .A2(\i_ibex/cs_registers_i/_0286_ ));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1420_  (.Y(\i_ibex/cs_registers_i/_0289_ ),
    .B(\i_ibex/cs_registers_i/_0160_ ),
    .A_N(\i_ibex/cs_registers_i/_0288_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1421_  (.Y(\i_ibex/cs_registers_i/_0290_ ),
    .B1(net450),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [2]),
    .A2(net988),
    .A1(net6),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1422_  (.B1(\i_ibex/cs_registers_i/_0290_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0291_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0285_ ),
    .A2(\i_ibex/cs_registers_i/_0289_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1423_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net466),
    .A2(\i_ibex/cs_registers_i/_0281_ ),
    .Y(\i_ibex/cs_registers_i/_0292_ ),
    .B1(\i_ibex/cs_registers_i/_0291_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1424_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net975),
    .Y(\i_ibex/csr_rdata [2]),
    .A2(\i_ibex/cs_registers_i/_0292_ ),
    .A1(\i_ibex/cs_registers_i/_0271_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1425_  (.Y(\i_ibex/cs_registers_i/_0293_ ),
    .A(net690),
    .B(\i_ibex/csr_rdata [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1426_  (.Y(\i_ibex/cs_registers_i/_0294_ ),
    .A(net541),
    .B(net631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1427_  (.B1(\i_ibex/cs_registers_i/_0294_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [2]),
    .VSS(VSS),
    .A1(net541),
    .A2(\i_ibex/cs_registers_i/_0293_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1428_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0295_ ),
    .A(net689),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1429_  (.A(net587),
    .B(\i_ibex/cs_registers_i/_0047_ ),
    .Y(\i_ibex/cs_registers_i/_0296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/_1430_  (.B(net589),
    .C(net7),
    .Y(\i_ibex/cs_registers_i/_0297_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net506));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1431_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0197_ ),
    .A2(\i_ibex/cs_registers_i/_0297_ ),
    .Y(\i_ibex/cs_registers_i/_0298_ ),
    .B1(net1065));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1432_  (.B1(\i_ibex/cs_registers_i/_0124_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0299_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0296_ ),
    .A2(\i_ibex/cs_registers_i/_0298_ ));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1433_  (.S0(net1063),
    .A0(\i_ibex/cs_registers_i/mscratch_q [1]),
    .A1(\i_ibex/csr_mepc [1]),
    .A2(\i_ibex/cs_registers_i/mcause_q [1]),
    .A3(\i_ibex/cs_registers_i/mtval_q [1]),
    .S1(net521),
    .X(\i_ibex/cs_registers_i/_0300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1434_  (.B(net453),
    .C(\i_ibex/cs_registers_i/_0300_ ),
    .A(net1061),
    .Y(\i_ibex/cs_registers_i/_0301_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1435_  (.A2(\i_ibex/cs_registers_i/_0301_ ),
    .A1(\i_ibex/cs_registers_i/_0299_ ),
    .B1(net1089),
    .X(\i_ibex/cs_registers_i/_0302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1436_  (.A(net519),
    .B_N(\i_ibex/cs_registers_i/mhpmcounter [2017]),
    .Y(\i_ibex/cs_registers_i/_0303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1437_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net519),
    .A2(\i_ibex/cs_registers_i/minstret_raw [33]),
    .Y(\i_ibex/cs_registers_i/_0304_ ),
    .B1(\i_ibex/cs_registers_i/_0303_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1438_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1985]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [1]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1439_  (.Y(\i_ibex/cs_registers_i/_0306_ ),
    .A(net463),
    .B(\i_ibex/cs_registers_i/_0305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1440_  (.B1(\i_ibex/cs_registers_i/_0306_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0307_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0243_ ),
    .A2(\i_ibex/cs_registers_i/_0304_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1441_  (.Y(\i_ibex/cs_registers_i/_0308_ ),
    .B1(\i_ibex/cs_registers_i/_0307_ ),
    .B2(\i_ibex/cs_registers_i/_0106_ ),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1442_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [1]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [1]),
    .A2(\i_ibex/csr_depc [1]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [1]),
    .S1(net1099),
    .X(\i_ibex/cs_registers_i/_0309_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1443_  (.Y(\i_ibex/cs_registers_i/_0310_ ),
    .B1(\i_ibex/cs_registers_i/_0309_ ),
    .B2(net461),
    .A2(net984),
    .A1(\i_ibex/csr_mtvec [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/cs_registers_i/_1444_  (.X(\i_ibex/cs_registers_i/_0311_ ),
    .A(\i_ibex/cs_registers_i/_0302_ ),
    .B(\i_ibex/cs_registers_i/_0308_ ),
    .C(\i_ibex/cs_registers_i/_0310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1445_  (.A(\i_ibex/cs_registers_i/_0295_ ),
    .B(net976),
    .C(\i_ibex/cs_registers_i/_0311_ ),
    .Y(\i_ibex/cs_registers_i/_0312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1446_  (.A0(\i_ibex/cs_registers_i/_0312_ ),
    .A1(net631),
    .S(net537),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1447_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2016]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [32]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1448_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [0]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0314_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1449_  (.Y(\i_ibex/cs_registers_i/_0315_ ),
    .B1(\i_ibex/cs_registers_i/_0314_ ),
    .B2(net462),
    .A2(\i_ibex/cs_registers_i/_0313_ ),
    .A1(\i_ibex/cs_registers_i/_0108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1450_  (.Y(\i_ibex/cs_registers_i/_0316_ ),
    .B(\i_ibex/cs_registers_i/_0106_ ),
    .A_N(\i_ibex/cs_registers_i/_0315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1451_  (.A(\i_ibex/cs_registers_i/mtval_q [0]),
    .B(net1063),
    .X(\i_ibex/cs_registers_i/_0317_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1452_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcause_q [0]),
    .A2(net1034),
    .Y(\i_ibex/cs_registers_i/_0318_ ),
    .B1(\i_ibex/cs_registers_i/_0317_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1453_  (.A(net1088),
    .B(\i_ibex/cs_registers_i/_0196_ ),
    .C(\i_ibex/cs_registers_i/_0197_ ),
    .D(\i_ibex/cs_registers_i/_0318_ ),
    .Y(\i_ibex/cs_registers_i/_0319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1454_  (.Y(\i_ibex/cs_registers_i/_0320_ ),
    .B1(\i_ibex/cs_registers_i/_0120_ ),
    .B2(\i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y [192]),
    .A2(net473),
    .A1(\i_ibex/cs_registers_i/mscratch_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1455_  (.A(\i_ibex/cs_registers_i/_0118_ ),
    .B(\i_ibex/cs_registers_i/_0320_ ),
    .Y(\i_ibex/cs_registers_i/_0321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1456_  (.B1(net465),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0322_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0319_ ),
    .A2(\i_ibex/cs_registers_i/_0321_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1457_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net8),
    .A2(\i_ibex/cs_registers_i/_0073_ ),
    .Y(\i_ibex/cs_registers_i/_0323_ ),
    .B1(\i_ibex/cs_registers_i/_0074_ ));
 sg13g2_inv_2 \i_ibex/cs_registers_i/_1458_  (.Y(\i_ibex/cs_registers_i/_0324_ ),
    .A(net1089),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1459_  (.Y(\i_ibex/cs_registers_i/_0325_ ),
    .A(net1035),
    .B(\i_ibex/cs_registers_i/_0324_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1460_  (.A(\i_ibex/cs_registers_i/_0323_ ),
    .B(\i_ibex/cs_registers_i/_0325_ ),
    .Y(\i_ibex/cs_registers_i/_0326_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1461_  (.Y(\i_ibex/cs_registers_i/_0327_ ),
    .B1(\i_ibex/cs_registers_i/_0124_ ),
    .B2(\i_ibex/cs_registers_i/_0326_ ),
    .A2(\i_ibex/cs_registers_i/_0082_ ),
    .A1(\i_ibex/csr_mepc [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1462_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [0]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [0]),
    .A2(\i_ibex/csr_depc [0]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [0]),
    .S1(net1100),
    .X(\i_ibex/cs_registers_i/_0328_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_2 \i_ibex/cs_registers_i/_1463_  (.A(net1094),
    .B(net1092),
    .C(\i_ibex/cs_registers_i/_0061_ ),
    .D(\i_ibex/cs_registers_i/_0062_ ),
    .X(\i_ibex/cs_registers_i/_0329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1464_  (.A(net519),
    .B_N(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_q ),
    .Y(\i_ibex/cs_registers_i/_0330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1465_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [0]),
    .A2(net519),
    .Y(\i_ibex/cs_registers_i/_0331_ ),
    .B1(\i_ibex/cs_registers_i/_0330_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1466_  (.A(net587),
    .B(\i_ibex/cs_registers_i/_0329_ ),
    .C(\i_ibex/cs_registers_i/_0325_ ),
    .D(\i_ibex/cs_registers_i/_0331_ ),
    .Y(\i_ibex/cs_registers_i/_0332_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1467_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net460),
    .C1(\i_ibex/cs_registers_i/_0332_ ),
    .B1(\i_ibex/cs_registers_i/_0328_ ),
    .A1(\i_ibex/csr_mtvec [0]),
    .Y(\i_ibex/cs_registers_i/_0333_ ),
    .A2(net984));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1468_  (.A(\i_ibex/cs_registers_i/_0316_ ),
    .B(\i_ibex/cs_registers_i/_0322_ ),
    .C(\i_ibex/cs_registers_i/_0327_ ),
    .D(\i_ibex/cs_registers_i/_0333_ ),
    .X(\i_ibex/cs_registers_i/_0334_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1469_  (.A(\i_ibex/cs_registers_i/_0295_ ),
    .B(net976),
    .C(\i_ibex/cs_registers_i/_0334_ ),
    .Y(\i_ibex/cs_registers_i/_0335_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1470_  (.A0(\i_ibex/cs_registers_i/_0335_ ),
    .A1(net631),
    .S(net1514),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1471_  (.A(\i_ibex/csr_mepc [30]),
    .B(net1069),
    .X(\i_ibex/cs_registers_i/_0336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1472_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [30]),
    .A2(net1039),
    .Y(\i_ibex/cs_registers_i/_0337_ ),
    .B1(\i_ibex/cs_registers_i/_0336_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1473_  (.B(net1072),
    .C(net508),
    .A(\i_ibex/cs_registers_i/mtval_q [30]),
    .Y(\i_ibex/cs_registers_i/_0338_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1474_  (.B1(\i_ibex/cs_registers_i/_0338_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0339_ ),
    .VSS(VSS),
    .A1(net511),
    .A2(\i_ibex/cs_registers_i/_0337_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1475_  (.Y(\i_ibex/cs_registers_i/_0340_ ),
    .B1(\i_ibex/cs_registers_i/_0339_ ),
    .B2(\i_ibex/cs_registers_i/_0025_ ),
    .A2(\i_ibex/cs_registers_i/_0087_ ),
    .A1(irqs_i[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout969 (.A(net970),
    .X(net969),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1477_  (.Y(\i_ibex/cs_registers_i/_0342_ ),
    .B(net454),
    .A_N(\i_ibex/cs_registers_i/_0340_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1478_  (.A(net1089),
    .B(\i_ibex/cs_registers_i/_0047_ ),
    .Y(\i_ibex/cs_registers_i/_0343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1479_  (.Y(\i_ibex/cs_registers_i/_0344_ ),
    .B1(net1031),
    .B2(\i_ibex/cs_registers_i/mie_q [14]),
    .A2(\i_ibex/cs_registers_i/_0343_ ),
    .A1(\i_ibex/csr_mtvec [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1480_  (.Y(\i_ibex/cs_registers_i/_0345_ ),
    .A(net589),
    .B(\i_ibex/cs_registers_i/_0115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1481_  (.B(\i_ibex/cs_registers_i/_0044_ ),
    .C(net462),
    .A(net465),
    .Y(\i_ibex/cs_registers_i/_0346_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1482_  (.B1(\i_ibex/cs_registers_i/_0346_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0347_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0344_ ),
    .A2(\i_ibex/cs_registers_i/_0345_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1483_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net9),
    .A2(net991),
    .Y(\i_ibex/cs_registers_i/_0348_ ),
    .B1(\i_ibex/cs_registers_i/_0347_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1484_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2014]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [30]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0349_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1485_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [30]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [30]),
    .A2(\i_ibex/csr_depc [30]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [30]),
    .S1(net1101),
    .X(\i_ibex/cs_registers_i/_0350_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1486_  (.Y(\i_ibex/cs_registers_i/_0351_ ),
    .B1(\i_ibex/cs_registers_i/_0350_ ),
    .B2(net461),
    .A2(\i_ibex/cs_registers_i/_0349_ ),
    .A1(net1004),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1487_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2046]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [62]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0352_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1488_  (.Y(\i_ibex/cs_registers_i/_0353_ ),
    .B1(net1002),
    .B2(\i_ibex/cs_registers_i/_0352_ ),
    .A2(net449),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1489_  (.A(\i_ibex/cs_registers_i/_0342_ ),
    .B(\i_ibex/cs_registers_i/_0348_ ),
    .C(\i_ibex/cs_registers_i/_0351_ ),
    .D(\i_ibex/cs_registers_i/_0353_ ),
    .X(\i_ibex/cs_registers_i/_0354_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1490_  (.A(\i_ibex/alu_operand_a_ex [30]),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0354_ ),
    .Y(\i_ibex/cs_registers_i/_0355_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/cs_registers_i/_1491_  (.A2(net633),
    .A1(\i_ibex/alu_operand_a_ex [30]),
    .B1(\i_ibex/cs_registers_i/_0355_ ),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1492_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2037]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [53]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0356_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1493_  (.A(net520),
    .B_N(\i_ibex/cs_registers_i/mhpmcounter [2005]),
    .Y(\i_ibex/cs_registers_i/_0357_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1494_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net520),
    .A2(\i_ibex/cs_registers_i/minstret_raw [21]),
    .Y(\i_ibex/cs_registers_i/_0358_ ),
    .B1(\i_ibex/cs_registers_i/_0357_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1495_  (.A(\i_ibex/cs_registers_i/_0218_ ),
    .B(\i_ibex/cs_registers_i/_0358_ ),
    .Y(\i_ibex/cs_registers_i/_0359_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1496_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0356_ ),
    .C1(\i_ibex/cs_registers_i/_0359_ ),
    .B1(net1002),
    .A1(net10),
    .Y(\i_ibex/cs_registers_i/_0360_ ),
    .A2(net990));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1497_  (.A0(\i_ibex/csr_mepc [21]),
    .A1(\i_ibex/cs_registers_i/mtval_q [21]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0361_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1498_  (.A(net589),
    .B_N(net1072),
    .Y(\i_ibex/cs_registers_i/_0362_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/cs_registers_i/_1499_  (.A(\i_ibex/cs_registers_i/_0324_ ),
    .B(\i_ibex/cs_registers_i/_0362_ ),
    .X(\i_ibex/cs_registers_i/_0363_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1500_  (.A0(\i_ibex/cs_registers_i/mscratch_q [21]),
    .A1(irqs_i[5]),
    .S(net587),
    .X(\i_ibex/cs_registers_i/_0364_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1501_  (.Y(\i_ibex/cs_registers_i/_0365_ ),
    .B1(\i_ibex/cs_registers_i/_0364_ ),
    .B2(net1031),
    .A2(\i_ibex/cs_registers_i/_0363_ ),
    .A1(\i_ibex/cs_registers_i/_0361_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1502_  (.A(\i_ibex/cs_registers_i/_0072_ ),
    .B(\i_ibex/cs_registers_i/_0365_ ),
    .Y(\i_ibex/cs_registers_i/_0366_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1503_  (.A0(\i_ibex/csr_mstatus_tw ),
    .A1(\i_ibex/cs_registers_i/mie_q [5]),
    .S(net587),
    .X(\i_ibex/cs_registers_i/_0367_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1504_  (.Y(\i_ibex/cs_registers_i/_0368_ ),
    .A(net1031),
    .B(\i_ibex/cs_registers_i/_0367_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1505_  (.B(net589),
    .C(\i_ibex/cs_registers_i/_0343_ ),
    .A(\i_ibex/csr_mtvec [21]),
    .Y(\i_ibex/cs_registers_i/_0369_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_1506_  (.Y(\i_ibex/cs_registers_i/_0370_ ),
    .A(net464),
    .B(\i_ibex/cs_registers_i/_0259_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1507_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0368_ ),
    .A2(\i_ibex/cs_registers_i/_0369_ ),
    .Y(\i_ibex/cs_registers_i/_0371_ ),
    .B1(\i_ibex/cs_registers_i/_0370_ ));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1508_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [21]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [21]),
    .A2(\i_ibex/csr_depc [21]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [21]),
    .S1(net1102),
    .X(\i_ibex/cs_registers_i/_0372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1509_  (.A(net459),
    .B(\i_ibex/cs_registers_i/_0372_ ),
    .X(\i_ibex/cs_registers_i/_0373_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1510_  (.A2(net447),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [21]),
    .B1(\i_ibex/cs_registers_i/_0373_ ),
    .X(\i_ibex/cs_registers_i/_0374_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1511_  (.A(net983),
    .B(\i_ibex/cs_registers_i/_0366_ ),
    .C(\i_ibex/cs_registers_i/_0371_ ),
    .D(\i_ibex/cs_registers_i/_0374_ ),
    .Y(\i_ibex/cs_registers_i/_0375_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1512_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net978),
    .Y(\i_ibex/csr_rdata [21]),
    .A2(\i_ibex/cs_registers_i/_0375_ ),
    .A1(\i_ibex/cs_registers_i/_0360_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1513_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net690),
    .A2(\i_ibex/csr_rdata [21]),
    .Y(\i_ibex/cs_registers_i/_0376_ ),
    .B1(net580));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1514_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0376_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [21]),
    .A2(\i_ibex/cs_registers_i/_0228_ ),
    .A1(net580));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1515_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2004]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [20]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0377_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1516_  (.Y(\i_ibex/cs_registers_i/_0378_ ),
    .B1(net1005),
    .B2(\i_ibex/cs_registers_i/_0377_ ),
    .A2(net449),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1517_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [52]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0379_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1518_  (.Y(\i_ibex/cs_registers_i/_0380_ ),
    .B1(net1000),
    .B2(\i_ibex/cs_registers_i/_0379_ ),
    .A2(net990),
    .A1(net11),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1519_  (.A0(\i_ibex/csr_mepc [20]),
    .A1(\i_ibex/cs_registers_i/mtval_q [20]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0381_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1520_  (.Y(\i_ibex/cs_registers_i/_0382_ ),
    .B1(\i_ibex/cs_registers_i/_0381_ ),
    .B2(net1070),
    .A2(net1040),
    .A1(\i_ibex/cs_registers_i/mscratch_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1521_  (.Y(\i_ibex/cs_registers_i/_0383_ ),
    .A(irqs_i[4]),
    .B(net457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1522_  (.B1(\i_ibex/cs_registers_i/_0383_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0384_ ),
    .VSS(VSS),
    .A1(net1033),
    .A2(\i_ibex/cs_registers_i/_0382_ ));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1523_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [20]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [20]),
    .A2(\i_ibex/csr_depc [20]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [20]),
    .S1(net1103),
    .X(\i_ibex/cs_registers_i/_0385_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1524_  (.Y(\i_ibex/cs_registers_i/_0386_ ),
    .B1(net1031),
    .B2(\i_ibex/cs_registers_i/mie_q [4]),
    .A2(\i_ibex/cs_registers_i/_0343_ ),
    .A1(\i_ibex/csr_mtvec [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1525_  (.B1(\i_ibex/cs_registers_i/_0346_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0387_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0345_ ),
    .A2(\i_ibex/cs_registers_i/_0386_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1526_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net461),
    .C1(\i_ibex/cs_registers_i/_0387_ ),
    .B1(\i_ibex/cs_registers_i/_0385_ ),
    .A1(net455),
    .Y(\i_ibex/cs_registers_i/_0388_ ),
    .A2(\i_ibex/cs_registers_i/_0384_ ));
 sg13g2_and3_2 \i_ibex/cs_registers_i/_1527_  (.X(\i_ibex/cs_registers_i/_0389_ ),
    .A(\i_ibex/cs_registers_i/_0378_ ),
    .B(\i_ibex/cs_registers_i/_0380_ ),
    .C(\i_ibex/cs_registers_i/_0388_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1528_  (.A(net578),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0389_ ),
    .Y(\i_ibex/cs_registers_i/_0390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/cs_registers_i/_1529_  (.A2(net633),
    .A1(net578),
    .B1(\i_ibex/cs_registers_i/_0390_ ),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout968 (.A(net970),
    .X(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout967 (.A(net970),
    .X(net967),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1533_  (.Y(\i_ibex/cs_registers_i/_0394_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [19]),
    .A2(net991),
    .A1(net12),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout965 (.A(net967),
    .X(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1535_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2035]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [51]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0396_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1536_  (.A(net1101),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [19]),
    .Y(\i_ibex/cs_registers_i/_0397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1537_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [19]),
    .A2(net1102),
    .Y(\i_ibex/cs_registers_i/_0398_ ),
    .B1(\i_ibex/cs_registers_i/_0397_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1538_  (.B(net1036),
    .C(net512),
    .A(\i_ibex/cs_registers_i/dscratch0_q [19]),
    .Y(\i_ibex/cs_registers_i/_0399_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1539_  (.B1(\i_ibex/cs_registers_i/_0399_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0400_ ),
    .VSS(VSS),
    .A1(net510),
    .A2(\i_ibex/cs_registers_i/_0398_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1540_  (.Y(\i_ibex/cs_registers_i/_0401_ ),
    .B1(\i_ibex/cs_registers_i/_0400_ ),
    .B2(net460),
    .A2(\i_ibex/cs_registers_i/_0396_ ),
    .A1(net1001),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1541_  (.A(\i_ibex/cs_registers_i/_0394_ ),
    .B(\i_ibex/cs_registers_i/_0401_ ),
    .X(\i_ibex/cs_registers_i/_0402_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1542_  (.A0(\i_ibex/csr_mepc [19]),
    .A1(\i_ibex/cs_registers_i/mtval_q [19]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0403_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1543_  (.Y(\i_ibex/cs_registers_i/_0404_ ),
    .B1(\i_ibex/cs_registers_i/_0403_ ),
    .B2(net1071),
    .A2(net1040),
    .A1(\i_ibex/cs_registers_i/mscratch_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1544_  (.Y(\i_ibex/cs_registers_i/_0405_ ),
    .A(irqs_i[3]),
    .B(net457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1545_  (.B1(\i_ibex/cs_registers_i/_0405_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0406_ ),
    .VSS(VSS),
    .A1(net1033),
    .A2(\i_ibex/cs_registers_i/_0404_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1546_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [19]),
    .C1(net983),
    .B1(net446),
    .A1(\i_ibex/cs_registers_i/mie_q [3]),
    .Y(\i_ibex/cs_registers_i/_0407_ ),
    .A2(net437));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1547_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [19]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0408_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1548_  (.Y(\i_ibex/cs_registers_i/_0409_ ),
    .B1(net1005),
    .B2(\i_ibex/cs_registers_i/_0408_ ),
    .A2(net986),
    .A1(\i_ibex/csr_mtvec [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1549_  (.Y(\i_ibex/cs_registers_i/_0410_ ),
    .A(\i_ibex/cs_registers_i/_0407_ ),
    .B(\i_ibex/cs_registers_i/_0409_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1550_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net454),
    .A2(\i_ibex/cs_registers_i/_0406_ ),
    .Y(\i_ibex/cs_registers_i/_0411_ ),
    .B1(\i_ibex/cs_registers_i/_0410_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1551_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net977),
    .Y(\i_ibex/csr_rdata [19]),
    .A2(\i_ibex/cs_registers_i/_0411_ ),
    .A1(\i_ibex/cs_registers_i/_0402_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1552_  (.Y(\i_ibex/cs_registers_i/_0412_ ),
    .A(net692),
    .B(\i_ibex/csr_rdata [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1553_  (.Y(\i_ibex/cs_registers_i/_0413_ ),
    .A(net576),
    .B(net631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1554_  (.B1(\i_ibex/cs_registers_i/_0413_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [19]),
    .VSS(VSS),
    .A1(net576),
    .A2(\i_ibex/cs_registers_i/_0412_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1555_  (.Y(\i_ibex/cs_registers_i/_0414_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [18]),
    .A2(net991),
    .A1(net13),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1556_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2034]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [50]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0415_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1557_  (.A(net1101),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [18]),
    .Y(\i_ibex/cs_registers_i/_0416_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1558_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [18]),
    .A2(net1101),
    .Y(\i_ibex/cs_registers_i/_0417_ ),
    .B1(\i_ibex/cs_registers_i/_0416_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1559_  (.B(net1036),
    .C(net512),
    .A(\i_ibex/cs_registers_i/dscratch0_q [18]),
    .Y(\i_ibex/cs_registers_i/_0418_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1560_  (.B1(\i_ibex/cs_registers_i/_0418_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0419_ ),
    .VSS(VSS),
    .A1(net510),
    .A2(\i_ibex/cs_registers_i/_0417_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1561_  (.Y(\i_ibex/cs_registers_i/_0420_ ),
    .B1(\i_ibex/cs_registers_i/_0419_ ),
    .B2(net460),
    .A2(\i_ibex/cs_registers_i/_0415_ ),
    .A1(net1001),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1562_  (.A(\i_ibex/cs_registers_i/_0414_ ),
    .B(\i_ibex/cs_registers_i/_0420_ ),
    .X(\i_ibex/cs_registers_i/_0421_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1563_  (.A0(\i_ibex/csr_mepc [18]),
    .A1(\i_ibex/cs_registers_i/mtval_q [18]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0422_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1564_  (.Y(\i_ibex/cs_registers_i/_0423_ ),
    .B1(\i_ibex/cs_registers_i/_0422_ ),
    .B2(net1071),
    .A2(net1040),
    .A1(\i_ibex/cs_registers_i/mscratch_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1565_  (.Y(\i_ibex/cs_registers_i/_0424_ ),
    .A(irqs_i[2]),
    .B(net457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1566_  (.B1(\i_ibex/cs_registers_i/_0424_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0425_ ),
    .VSS(VSS),
    .A1(net1033),
    .A2(\i_ibex/cs_registers_i/_0423_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1567_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [18]),
    .C1(net982),
    .B1(net446),
    .A1(\i_ibex/cs_registers_i/mie_q [2]),
    .Y(\i_ibex/cs_registers_i/_0426_ ),
    .A2(net437));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1568_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2002]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [18]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0427_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1569_  (.Y(\i_ibex/cs_registers_i/_0428_ ),
    .B1(net1005),
    .B2(\i_ibex/cs_registers_i/_0427_ ),
    .A2(net985),
    .A1(\i_ibex/csr_mtvec [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1570_  (.Y(\i_ibex/cs_registers_i/_0429_ ),
    .A(\i_ibex/cs_registers_i/_0426_ ),
    .B(\i_ibex/cs_registers_i/_0428_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1571_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net454),
    .A2(\i_ibex/cs_registers_i/_0425_ ),
    .Y(\i_ibex/cs_registers_i/_0430_ ),
    .B1(\i_ibex/cs_registers_i/_0429_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1572_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net977),
    .Y(\i_ibex/csr_rdata [18]),
    .A2(\i_ibex/cs_registers_i/_0430_ ),
    .A1(\i_ibex/cs_registers_i/_0421_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1573_  (.Y(\i_ibex/cs_registers_i/_0431_ ),
    .A(net692),
    .B(\i_ibex/csr_rdata [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1574_  (.Y(\i_ibex/cs_registers_i/_0432_ ),
    .A(net574),
    .B(net631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1575_  (.B1(\i_ibex/cs_registers_i/_0432_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [18]),
    .VSS(VSS),
    .A1(net574),
    .A2(\i_ibex/cs_registers_i/_0431_ ));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1576_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [17]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [17]),
    .A2(\i_ibex/csr_depc [17]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [17]),
    .S1(net1101),
    .X(\i_ibex/cs_registers_i/_0433_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1577_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2001]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [17]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0434_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1578_  (.Y(\i_ibex/cs_registers_i/_0435_ ),
    .B1(\i_ibex/cs_registers_i/_0434_ ),
    .B2(net1005),
    .A2(\i_ibex/cs_registers_i/_0433_ ),
    .A1(net459),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1579_  (.Y(\i_ibex/cs_registers_i/_0436_ ),
    .B1(net991),
    .B2(net14),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1580_  (.A(\i_ibex/cs_registers_i/_0435_ ),
    .B(\i_ibex/cs_registers_i/_0436_ ),
    .X(\i_ibex/cs_registers_i/_0437_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1581_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2033]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [49]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0438_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1582_  (.A0(\i_ibex/cs_registers_i/mscratch_q [17]),
    .A1(irqs_i[1]),
    .S(net587),
    .X(\i_ibex/cs_registers_i/_0439_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1583_  (.A0(\i_ibex/csr_mepc [17]),
    .A1(\i_ibex/cs_registers_i/mtval_q [17]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0440_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1584_  (.Y(\i_ibex/cs_registers_i/_0441_ ),
    .B1(\i_ibex/cs_registers_i/_0440_ ),
    .B2(\i_ibex/cs_registers_i/_0363_ ),
    .A2(\i_ibex/cs_registers_i/_0439_ ),
    .A1(\i_ibex/cs_registers_i/_0086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1585_  (.Y(\i_ibex/cs_registers_i/_0442_ ),
    .B(\i_ibex/cs_registers_i/_0120_ ),
    .A_N(\i_ibex/cs_registers_i/_0118_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1586_  (.B1(\i_ibex/cs_registers_i/_0442_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0443_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0196_ ),
    .A2(\i_ibex/cs_registers_i/_0441_ ));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1587_  (.Y(\i_ibex/cs_registers_i/_0444_ ),
    .B(\i_ibex/cs_registers_i/mstatus_q [1]),
    .A_N(net1066),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1588_  (.B(net1072),
    .C(net587),
    .A(\i_ibex/csr_mtvec [17]),
    .Y(\i_ibex/cs_registers_i/_0445_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1589_  (.B1(\i_ibex/cs_registers_i/_0445_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0446_ ),
    .VSS(VSS),
    .A1(net587),
    .A2(\i_ibex/cs_registers_i/_0444_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1590_  (.Y(\i_ibex/cs_registers_i/_0447_ ),
    .B1(\i_ibex/cs_registers_i/_0234_ ),
    .B2(\i_ibex/cs_registers_i/_0446_ ),
    .A2(net456),
    .A1(\i_ibex/cs_registers_i/mie_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1591_  (.A(\i_ibex/cs_registers_i/_0370_ ),
    .B(\i_ibex/cs_registers_i/_0447_ ),
    .Y(\i_ibex/cs_registers_i/_0448_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1592_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net464),
    .C1(\i_ibex/cs_registers_i/_0448_ ),
    .B1(\i_ibex/cs_registers_i/_0443_ ),
    .A1(net1002),
    .Y(\i_ibex/cs_registers_i/_0449_ ),
    .A2(\i_ibex/cs_registers_i/_0438_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1593_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net978),
    .Y(\i_ibex/csr_rdata [17]),
    .A2(\i_ibex/cs_registers_i/_0449_ ),
    .A1(\i_ibex/cs_registers_i/_0437_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1594_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net690),
    .A2(\i_ibex/csr_rdata [17]),
    .Y(\i_ibex/cs_registers_i/_0450_ ),
    .B1(net572));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1595_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0450_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [17]),
    .A2(\i_ibex/cs_registers_i/_0228_ ),
    .A1(net572));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1596_  (.Y(\i_ibex/cs_registers_i/_0451_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [16]),
    .A2(net990),
    .A1(net15),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1597_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2032]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [48]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0452_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1598_  (.A(net1101),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [16]),
    .Y(\i_ibex/cs_registers_i/_0453_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1599_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [16]),
    .A2(net1101),
    .Y(\i_ibex/cs_registers_i/_0454_ ),
    .B1(\i_ibex/cs_registers_i/_0453_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1600_  (.B(net1036),
    .C(net512),
    .A(\i_ibex/cs_registers_i/dscratch0_q [16]),
    .Y(\i_ibex/cs_registers_i/_0455_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1601_  (.B1(\i_ibex/cs_registers_i/_0455_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0456_ ),
    .VSS(VSS),
    .A1(net510),
    .A2(\i_ibex/cs_registers_i/_0454_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1602_  (.Y(\i_ibex/cs_registers_i/_0457_ ),
    .B1(\i_ibex/cs_registers_i/_0456_ ),
    .B2(net460),
    .A2(\i_ibex/cs_registers_i/_0452_ ),
    .A1(net1000),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1603_  (.A(\i_ibex/cs_registers_i/_0451_ ),
    .B(\i_ibex/cs_registers_i/_0457_ ),
    .X(\i_ibex/cs_registers_i/_0458_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1604_  (.A0(\i_ibex/csr_mepc [16]),
    .A1(\i_ibex/cs_registers_i/mtval_q [16]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0459_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1605_  (.Y(\i_ibex/cs_registers_i/_0460_ ),
    .B1(\i_ibex/cs_registers_i/_0459_ ),
    .B2(net1070),
    .A2(\i_ibex/cs_registers_i/_0026_ ),
    .A1(\i_ibex/cs_registers_i/mscratch_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1606_  (.Y(\i_ibex/cs_registers_i/_0461_ ),
    .A(irqs_i[0]),
    .B(net457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1607_  (.B1(\i_ibex/cs_registers_i/_0461_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0462_ ),
    .VSS(VSS),
    .A1(net1033),
    .A2(\i_ibex/cs_registers_i/_0460_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1608_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [16]),
    .C1(net982),
    .B1(net446),
    .A1(\i_ibex/cs_registers_i/mie_q [0]),
    .Y(\i_ibex/cs_registers_i/_0463_ ),
    .A2(net437));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1609_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2000]),
    .A1(net1494),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0464_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1610_  (.Y(\i_ibex/cs_registers_i/_0465_ ),
    .B1(net1004),
    .B2(\i_ibex/cs_registers_i/_0464_ ),
    .A2(net985),
    .A1(\i_ibex/csr_mtvec [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1611_  (.Y(\i_ibex/cs_registers_i/_0466_ ),
    .A(\i_ibex/cs_registers_i/_0463_ ),
    .B(\i_ibex/cs_registers_i/_0465_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1612_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net454),
    .A2(\i_ibex/cs_registers_i/_0462_ ),
    .Y(\i_ibex/cs_registers_i/_0467_ ),
    .B1(\i_ibex/cs_registers_i/_0466_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1613_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net977),
    .Y(\i_ibex/csr_rdata [16]),
    .A2(\i_ibex/cs_registers_i/_0467_ ),
    .A1(\i_ibex/cs_registers_i/_0458_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1614_  (.Y(\i_ibex/cs_registers_i/_0468_ ),
    .A(net691),
    .B(\i_ibex/csr_rdata [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1615_  (.Y(\i_ibex/cs_registers_i/_0469_ ),
    .A(net570),
    .B(net634),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1616_  (.B1(\i_ibex/cs_registers_i/_0469_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [16]),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_a_ex [16]),
    .A2(\i_ibex/cs_registers_i/_0468_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1617_  (.Y(\i_ibex/cs_registers_i/_0470_ ),
    .B1(net986),
    .B2(\i_ibex/csr_mtvec [15]),
    .A2(\i_ibex/cs_registers_i/_0082_ ),
    .A1(\i_ibex/csr_mepc [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1618_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2031]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [47]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0471_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout964 (.A(\i_ibex/cs_registers_i/csr_wdata_int [30]),
    .X(net964),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1620_  (.Y(\i_ibex/cs_registers_i/_0473_ ),
    .A(\i_ibex/cs_registers_i/mscratch_q [15]),
    .B(net1034),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1621_  (.B(net1062),
    .C(net508),
    .A(\i_ibex/cs_registers_i/mtval_q [15]),
    .Y(\i_ibex/cs_registers_i/_0474_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1622_  (.B1(\i_ibex/cs_registers_i/_0474_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0475_ ),
    .VSS(VSS),
    .A1(net507),
    .A2(\i_ibex/cs_registers_i/_0473_ ));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1623_  (.A(\i_ibex/cs_registers_i/_0118_ ),
    .B(\i_ibex/cs_registers_i/_0164_ ),
    .Y(\i_ibex/cs_registers_i/_0476_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1624_  (.A2(\i_ibex/cs_registers_i/_0475_ ),
    .A1(\i_ibex/cs_registers_i/_0272_ ),
    .B1(\i_ibex/cs_registers_i/_0476_ ),
    .X(\i_ibex/cs_registers_i/_0477_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1625_  (.Y(\i_ibex/cs_registers_i/_0478_ ),
    .B1(\i_ibex/cs_registers_i/_0477_ ),
    .B2(net466),
    .A2(\i_ibex/cs_registers_i/_0471_ ),
    .A1(net998),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1626_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [15]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0479_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1627_  (.Y(\i_ibex/cs_registers_i/_0480_ ),
    .B1(net1005),
    .B2(\i_ibex/cs_registers_i/_0479_ ),
    .A2(net990),
    .A1(net16),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1628_  (.A(net1100),
    .B_N(\i_ibex/debug_ebreakm ),
    .Y(\i_ibex/cs_registers_i/_0481_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1629_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0481_ ),
    .Y(\i_ibex/cs_registers_i/_0482_ ),
    .A2(net1105),
    .A1(\i_ibex/csr_depc [15]));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1630_  (.B(net1038),
    .C(net508),
    .A(\i_ibex/cs_registers_i/dscratch0_q [15]),
    .Y(\i_ibex/cs_registers_i/_0483_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1631_  (.B1(\i_ibex/cs_registers_i/_0483_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0484_ ),
    .VSS(VSS),
    .A1(net511),
    .A2(\i_ibex/cs_registers_i/_0482_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1632_  (.A(net459),
    .B(\i_ibex/cs_registers_i/_0484_ ),
    .X(\i_ibex/cs_registers_i/_0485_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1633_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [15]),
    .C1(\i_ibex/cs_registers_i/_0485_ ),
    .B1(net450),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [15]),
    .Y(\i_ibex/cs_registers_i/_0486_ ),
    .A2(net446));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1634_  (.A(\i_ibex/cs_registers_i/_0470_ ),
    .B(\i_ibex/cs_registers_i/_0478_ ),
    .C(\i_ibex/cs_registers_i/_0480_ ),
    .D(\i_ibex/cs_registers_i/_0486_ ),
    .X(\i_ibex/cs_registers_i/_0487_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1635_  (.A(\i_ibex/alu_operand_a_ex [15]),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0487_ ),
    .Y(\i_ibex/cs_registers_i/_0488_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/cs_registers_i/_1636_  (.A2(net633),
    .A1(\i_ibex/alu_operand_a_ex [15]),
    .B1(\i_ibex/cs_registers_i/_0488_ ),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1637_  (.Y(\i_ibex/cs_registers_i/_0489_ ),
    .A(\i_ibex/cs_registers_i/mscratch_q [14]),
    .B(net1034),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1638_  (.B(net1062),
    .C(net511),
    .A(\i_ibex/cs_registers_i/mtval_q [14]),
    .Y(\i_ibex/cs_registers_i/_0490_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1639_  (.B1(\i_ibex/cs_registers_i/_0490_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0491_ ),
    .VSS(VSS),
    .A1(net508),
    .A2(\i_ibex/cs_registers_i/_0489_ ));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1640_  (.A2(\i_ibex/cs_registers_i/_0491_ ),
    .A1(\i_ibex/cs_registers_i/_0272_ ),
    .B1(\i_ibex/cs_registers_i/_0476_ ),
    .X(\i_ibex/cs_registers_i/_0492_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1641_  (.Y(\i_ibex/cs_registers_i/_0493_ ),
    .B1(\i_ibex/cs_registers_i/_0492_ ),
    .B2(net466),
    .A2(\i_ibex/cs_registers_i/_0082_ ),
    .A1(\i_ibex/csr_mepc [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1642_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2030]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [46]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0494_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1643_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1998]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [14]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0495_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1644_  (.Y(\i_ibex/cs_registers_i/_0496_ ),
    .B1(\i_ibex/cs_registers_i/_0495_ ),
    .B2(net1003),
    .A2(\i_ibex/cs_registers_i/_0494_ ),
    .A1(net999),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1645_  (.Y(\i_ibex/cs_registers_i/_0497_ ),
    .B1(net989),
    .B2(net17),
    .A2(net449),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1646_  (.A(net1099),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [14]),
    .Y(\i_ibex/cs_registers_i/_0498_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1647_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [14]),
    .A2(net1099),
    .Y(\i_ibex/cs_registers_i/_0499_ ),
    .B1(\i_ibex/cs_registers_i/_0498_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1648_  (.B(\i_ibex/cs_registers_i/_0054_ ),
    .C(net510),
    .A(\i_ibex/cs_registers_i/dscratch0_q [14]),
    .Y(\i_ibex/cs_registers_i/_0500_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1649_  (.B1(\i_ibex/cs_registers_i/_0500_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0501_ ),
    .VSS(VSS),
    .A1(net507),
    .A2(\i_ibex/cs_registers_i/_0499_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1650_  (.A(net459),
    .B(\i_ibex/cs_registers_i/_0501_ ),
    .X(\i_ibex/cs_registers_i/_0502_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1651_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [14]),
    .C1(\i_ibex/cs_registers_i/_0502_ ),
    .B1(net450),
    .A1(\i_ibex/csr_mtvec [14]),
    .Y(\i_ibex/cs_registers_i/_0503_ ),
    .A2(net984));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1652_  (.A(\i_ibex/cs_registers_i/_0493_ ),
    .B(\i_ibex/cs_registers_i/_0496_ ),
    .C(\i_ibex/cs_registers_i/_0497_ ),
    .D(\i_ibex/cs_registers_i/_0503_ ),
    .X(\i_ibex/cs_registers_i/_0504_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1653_  (.A(net568),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0504_ ),
    .Y(\i_ibex/cs_registers_i/_0505_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1654_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0505_ ),
    .Y(\i_ibex/cs_registers_i/_0506_ ),
    .A2(net633),
    .A1(net568));
 sg13g2_inv_2 \i_ibex/cs_registers_i/_1655_  (.Y(\i_ibex/cs_registers_i/csr_wdata_int [14]),
    .A(\i_ibex/cs_registers_i/_0506_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1656_  (.Y(\i_ibex/cs_registers_i/_0507_ ),
    .B1(net987),
    .B2(\i_ibex/csr_mtvec [13]),
    .A2(\i_ibex/cs_registers_i/_0082_ ),
    .A1(\i_ibex/csr_mepc [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1657_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2029]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [45]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0508_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1658_  (.Y(\i_ibex/cs_registers_i/_0509_ ),
    .A(\i_ibex/cs_registers_i/mscratch_q [13]),
    .B(net1034),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1659_  (.B(net1062),
    .C(net508),
    .A(\i_ibex/cs_registers_i/mtval_q [13]),
    .Y(\i_ibex/cs_registers_i/_0510_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1660_  (.B1(\i_ibex/cs_registers_i/_0510_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0511_ ),
    .VSS(VSS),
    .A1(net511),
    .A2(\i_ibex/cs_registers_i/_0509_ ));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1661_  (.A2(\i_ibex/cs_registers_i/_0511_ ),
    .A1(\i_ibex/cs_registers_i/_0272_ ),
    .B1(\i_ibex/cs_registers_i/_0476_ ),
    .X(\i_ibex/cs_registers_i/_0512_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1662_  (.Y(\i_ibex/cs_registers_i/_0513_ ),
    .B1(\i_ibex/cs_registers_i/_0512_ ),
    .B2(net465),
    .A2(\i_ibex/cs_registers_i/_0508_ ),
    .A1(net998),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1663_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1997]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [13]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0514_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1664_  (.Y(\i_ibex/cs_registers_i/_0515_ ),
    .B1(net1003),
    .B2(\i_ibex/cs_registers_i/_0514_ ),
    .A2(net988),
    .A1(net18),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1665_  (.A(net1104),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [13]),
    .Y(\i_ibex/cs_registers_i/_0516_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1666_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [13]),
    .A2(net1104),
    .Y(\i_ibex/cs_registers_i/_0517_ ),
    .B1(\i_ibex/cs_registers_i/_0516_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1667_  (.B(net1038),
    .C(net508),
    .A(\i_ibex/cs_registers_i/dscratch0_q [13]),
    .Y(\i_ibex/cs_registers_i/_0518_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1668_  (.B1(\i_ibex/cs_registers_i/_0518_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0519_ ),
    .VSS(VSS),
    .A1(net511),
    .A2(\i_ibex/cs_registers_i/_0517_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1669_  (.A(net459),
    .B(\i_ibex/cs_registers_i/_0519_ ),
    .X(\i_ibex/cs_registers_i/_0520_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1670_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [13]),
    .C1(\i_ibex/cs_registers_i/_0520_ ),
    .B1(net450),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [13]),
    .Y(\i_ibex/cs_registers_i/_0521_ ),
    .A2(net446));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1671_  (.A(\i_ibex/cs_registers_i/_0507_ ),
    .B(\i_ibex/cs_registers_i/_0513_ ),
    .C(\i_ibex/cs_registers_i/_0515_ ),
    .D(\i_ibex/cs_registers_i/_0521_ ),
    .X(\i_ibex/cs_registers_i/_0522_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1672_  (.A(net566),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0522_ ),
    .Y(\i_ibex/cs_registers_i/_0523_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1673_  (.A2(net633),
    .A1(net566),
    .B1(\i_ibex/cs_registers_i/_0523_ ),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1674_  (.Y(\i_ibex/cs_registers_i/_0524_ ),
    .B(\i_ibex/cs_registers_i/mscratch_q [12]),
    .A_N(net507),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1675_  (.B(net1062),
    .C(net511),
    .A(\i_ibex/cs_registers_i/mtval_q [12]),
    .Y(\i_ibex/cs_registers_i/_0525_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1676_  (.B1(\i_ibex/cs_registers_i/_0525_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0526_ ),
    .VSS(VSS),
    .A1(net1064),
    .A2(\i_ibex/cs_registers_i/_0524_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1677_  (.A(\i_ibex/cs_registers_i/_0042_ ),
    .B(\i_ibex/cs_registers_i/_0256_ ),
    .Y(\i_ibex/cs_registers_i/_0527_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1678_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0527_ ),
    .C1(\i_ibex/cs_registers_i/_0254_ ),
    .B1(\i_ibex/cs_registers_i/_0526_ ),
    .A1(net19),
    .Y(\i_ibex/cs_registers_i/_0528_ ),
    .A2(net988));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1679_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [12]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0529_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1680_  (.A(net1066),
    .B(net589),
    .Y(\i_ibex/cs_registers_i/_0530_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1681_  (.A(net1034),
    .B(net1061),
    .Y(\i_ibex/cs_registers_i/_0531_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1682_  (.Y(\i_ibex/cs_registers_i/_0532_ ),
    .B1(\i_ibex/cs_registers_i/_0531_ ),
    .B2(\i_ibex/csr_mtvec [12]),
    .A2(\i_ibex/cs_registers_i/_0530_ ),
    .A1(\i_ibex/cs_registers_i/mstatus_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1683_  (.Y(\i_ibex/cs_registers_i/_0533_ ),
    .A(\i_ibex/cs_registers_i/_0259_ ),
    .B(\i_ibex/cs_registers_i/_0234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1684_  (.B(\i_ibex/cs_registers_i/_0286_ ),
    .C(net473),
    .A(\i_ibex/csr_mepc [12]),
    .Y(\i_ibex/cs_registers_i/_0534_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0071_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1685_  (.B1(\i_ibex/cs_registers_i/_0534_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0535_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0532_ ),
    .A2(\i_ibex/cs_registers_i/_0533_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1686_  (.Y(\i_ibex/cs_registers_i/_0536_ ),
    .B1(\i_ibex/cs_registers_i/_0535_ ),
    .B2(net464),
    .A2(\i_ibex/cs_registers_i/_0529_ ),
    .A1(net1003),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1687_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2028]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [44]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0537_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1688_  (.A(net1099),
    .B_N(\i_ibex/debug_ebreaku ),
    .Y(\i_ibex/cs_registers_i/_0538_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1689_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0538_ ),
    .Y(\i_ibex/cs_registers_i/_0539_ ),
    .A2(net1100),
    .A1(\i_ibex/csr_depc [12]));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1690_  (.B(net1068),
    .C(net509),
    .A(\i_ibex/cs_registers_i/dscratch1_q [12]),
    .Y(\i_ibex/cs_registers_i/_0540_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1691_  (.B1(\i_ibex/cs_registers_i/_0540_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0541_ ),
    .VSS(VSS),
    .A1(net508),
    .A2(\i_ibex/cs_registers_i/_0539_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1692_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [12]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [12]),
    .S(net1090),
    .X(\i_ibex/cs_registers_i/_0542_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/_1693_  (.X(\i_ibex/cs_registers_i/_0543_ ),
    .A(\i_ibex/cs_registers_i/_0135_ ),
    .B(\i_ibex/cs_registers_i/_0160_ ),
    .C(\i_ibex/cs_registers_i/_0542_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1694_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net460),
    .C1(\i_ibex/cs_registers_i/_0543_ ),
    .B1(\i_ibex/cs_registers_i/_0541_ ),
    .A1(net998),
    .Y(\i_ibex/cs_registers_i/_0544_ ),
    .A2(\i_ibex/cs_registers_i/_0537_ ));
 sg13g2_and3_1 \i_ibex/cs_registers_i/_1695_  (.X(\i_ibex/cs_registers_i/_0545_ ),
    .A(\i_ibex/cs_registers_i/_0528_ ),
    .B(\i_ibex/cs_registers_i/_0536_ ),
    .C(\i_ibex/cs_registers_i/_0544_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 \i_ibex/cs_registers_i/_1696_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0546_ ),
    .B(\i_ibex/cs_registers_i/_0545_ ),
    .A(net975));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1697_  (.A(net564),
    .B(\i_ibex/cs_registers_i/_0295_ ),
    .C(\i_ibex/cs_registers_i/_0546_ ),
    .Y(\i_ibex/cs_registers_i/_0547_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1698_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0547_ ),
    .Y(\i_ibex/cs_registers_i/_0548_ ),
    .A2(net633),
    .A1(net564));
 sg13g2_inv_2 \i_ibex/cs_registers_i/_1699_  (.Y(\i_ibex/cs_registers_i/csr_wdata_int [12]),
    .A(\i_ibex/cs_registers_i/_0548_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1700_  (.A(net520),
    .B_N(\i_ibex/cs_registers_i/mhpmcounter [2013]),
    .Y(\i_ibex/cs_registers_i/_0549_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1701_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net520),
    .A2(\i_ibex/cs_registers_i/minstret_raw [29]),
    .Y(\i_ibex/cs_registers_i/_0550_ ),
    .B1(\i_ibex/cs_registers_i/_0549_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1702_  (.A(\i_ibex/cs_registers_i/_0218_ ),
    .B(\i_ibex/cs_registers_i/_0550_ ),
    .Y(\i_ibex/cs_registers_i/_0551_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1703_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/dcsr_q [29]),
    .C1(\i_ibex/cs_registers_i/_0551_ ),
    .B1(net445),
    .A1(\i_ibex/csr_mtvec [29]),
    .Y(\i_ibex/cs_registers_i/_0552_ ),
    .A2(net987));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1704_  (.B(\i_ibex/cs_registers_i/_0059_ ),
    .C(net457),
    .A(net20),
    .Y(\i_ibex/cs_registers_i/_0553_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1705_  (.A(net1094),
    .B(\i_ibex/cs_registers_i/_0062_ ),
    .Y(\i_ibex/cs_registers_i/_0554_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1706_  (.Y(\i_ibex/cs_registers_i/_0555_ ),
    .A(\i_ibex/csr_depc [29]),
    .B(net1072),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/_1707_  (.B(net519),
    .C(\i_ibex/cs_registers_i/dscratch0_q [29]),
    .Y(\i_ibex/cs_registers_i/_0556_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1068));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1708_  (.B1(\i_ibex/cs_registers_i/_0556_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0557_ ),
    .VSS(VSS),
    .A1(net512),
    .A2(\i_ibex/cs_registers_i/_0555_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1709_  (.B(\i_ibex/cs_registers_i/_0554_ ),
    .C(\i_ibex/cs_registers_i/_0557_ ),
    .A(net1042),
    .Y(\i_ibex/cs_registers_i/_0558_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1710_  (.A2(\i_ibex/cs_registers_i/_0558_ ),
    .A1(\i_ibex/cs_registers_i/_0553_ ),
    .B1(\i_ibex/cs_registers_i/_0056_ ),
    .X(\i_ibex/cs_registers_i/_0559_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1711_  (.Y(\i_ibex/cs_registers_i/_0560_ ),
    .B1(net453),
    .B2(\i_ibex/cs_registers_i/mtval_q [29]),
    .A2(\i_ibex/cs_registers_i/_0127_ ),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1712_  (.Y(\i_ibex/cs_registers_i/_0561_ ),
    .B(\i_ibex/cs_registers_i/_0128_ ),
    .A_N(\i_ibex/cs_registers_i/_0560_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1713_  (.A(irqs_i[13]),
    .B(net589),
    .X(\i_ibex/cs_registers_i/_0562_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1714_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [29]),
    .A2(\i_ibex/cs_registers_i/_0013_ ),
    .Y(\i_ibex/cs_registers_i/_0563_ ),
    .B1(\i_ibex/cs_registers_i/_0562_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1715_  (.Y(\i_ibex/cs_registers_i/_0564_ ),
    .A(\i_ibex/csr_mepc [29]),
    .B(\i_ibex/cs_registers_i/_0362_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1716_  (.B1(\i_ibex/cs_registers_i/_0564_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0565_ ),
    .VSS(VSS),
    .A1(net1072),
    .A2(\i_ibex/cs_registers_i/_0563_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1717_  (.A(net453),
    .B(\i_ibex/cs_registers_i/_0234_ ),
    .X(\i_ibex/cs_registers_i/_0566_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1718_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0566_ ),
    .C1(\i_ibex/cs_registers_i/_0254_ ),
    .B1(\i_ibex/cs_registers_i/_0565_ ),
    .A1(\i_ibex/cs_registers_i/mie_q [13]),
    .Y(\i_ibex/cs_registers_i/_0567_ ),
    .A2(net436));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1719_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2045]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [61]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0568_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1720_  (.Y(\i_ibex/cs_registers_i/_0569_ ),
    .B1(net1002),
    .B2(\i_ibex/cs_registers_i/_0568_ ),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/_1721_  (.A(\i_ibex/cs_registers_i/_0559_ ),
    .B(\i_ibex/cs_registers_i/_0561_ ),
    .C(\i_ibex/cs_registers_i/_0567_ ),
    .D(\i_ibex/cs_registers_i/_0569_ ),
    .X(\i_ibex/cs_registers_i/_0570_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1722_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net975),
    .Y(\i_ibex/csr_rdata [29]),
    .A2(\i_ibex/cs_registers_i/_0570_ ),
    .A1(\i_ibex/cs_registers_i/_0552_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1723_  (.Y(\i_ibex/cs_registers_i/_0571_ ),
    .A(net690),
    .B(\i_ibex/csr_rdata [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1724_  (.Y(\i_ibex/cs_registers_i/_0572_ ),
    .A(\i_ibex/alu_operand_a_ex [29]),
    .B(net631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1725_  (.B1(\i_ibex/cs_registers_i/_0572_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [29]),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_a_ex [29]),
    .A2(\i_ibex/cs_registers_i/_0571_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1726_  (.A(net1099),
    .B_N(net507),
    .Y(\i_ibex/cs_registers_i/_0573_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1727_  (.A0(\i_ibex/csr_depc [11]),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [11]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0574_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1728_  (.Y(\i_ibex/cs_registers_i/_0575_ ),
    .B1(\i_ibex/cs_registers_i/_0574_ ),
    .B2(net1068),
    .A2(\i_ibex/cs_registers_i/_0573_ ),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1729_  (.A(\i_ibex/cs_registers_i/_0575_ ),
    .B_N(net461),
    .Y(\i_ibex/cs_registers_i/_0576_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1730_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net21),
    .C1(\i_ibex/cs_registers_i/_0576_ ),
    .B1(net989),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [11]),
    .Y(\i_ibex/cs_registers_i/_0577_ ),
    .A2(net449));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1731_  (.A0(\i_ibex/csr_mepc [11]),
    .A1(\i_ibex/cs_registers_i/mtval_q [11]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0578_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1732_  (.A0(\i_ibex/cs_registers_i/mscratch_q [11]),
    .A1(net22),
    .S(net587),
    .X(\i_ibex/cs_registers_i/_0579_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1733_  (.Y(\i_ibex/cs_registers_i/_0580_ ),
    .B1(\i_ibex/cs_registers_i/_0579_ ),
    .B2(net1031),
    .A2(\i_ibex/cs_registers_i/_0578_ ),
    .A1(\i_ibex/cs_registers_i/_0363_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1734_  (.B1(\i_ibex/cs_registers_i/_0442_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0581_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0196_ ),
    .A2(\i_ibex/cs_registers_i/_0580_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1735_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0582_ ),
    .A(\i_ibex/cs_registers_i/_0106_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1736_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1995]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [11]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0583_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1737_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2027]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [43]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0584_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1738_  (.Y(\i_ibex/cs_registers_i/_0585_ ),
    .B1(\i_ibex/cs_registers_i/_0584_ ),
    .B2(\i_ibex/cs_registers_i/_0108_ ),
    .A2(\i_ibex/cs_registers_i/_0583_ ),
    .A1(net462),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1739_  (.A0(\i_ibex/cs_registers_i/mie_q [16]),
    .A1(\i_ibex/csr_mtvec [11]),
    .S(net1072),
    .X(\i_ibex/cs_registers_i/_0586_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1740_  (.A(net1100),
    .B_N(\i_ibex/cs_registers_i/mstatus_q [2]),
    .Y(\i_ibex/cs_registers_i/_0587_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1741_  (.A0(\i_ibex/cs_registers_i/_0586_ ),
    .A1(\i_ibex/cs_registers_i/_0587_ ),
    .S(net1061),
    .X(\i_ibex/cs_registers_i/_0588_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1742_  (.B(\i_ibex/cs_registers_i/_0234_ ),
    .C(\i_ibex/cs_registers_i/_0588_ ),
    .A(\i_ibex/cs_registers_i/_0115_ ),
    .Y(\i_ibex/cs_registers_i/_0589_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1743_  (.B1(\i_ibex/cs_registers_i/_0589_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0590_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0582_ ),
    .A2(\i_ibex/cs_registers_i/_0585_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1744_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net464),
    .C1(\i_ibex/cs_registers_i/_0590_ ),
    .B1(\i_ibex/cs_registers_i/_0581_ ),
    .A1(\i_ibex/cs_registers_i/dcsr_q [11]),
    .Y(\i_ibex/cs_registers_i/_0591_ ),
    .A2(\i_ibex/cs_registers_i/_0161_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1745_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net975),
    .Y(\i_ibex/csr_rdata [11]),
    .A2(\i_ibex/cs_registers_i/_0591_ ),
    .A1(\i_ibex/cs_registers_i/_0577_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1746_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net691),
    .A2(\i_ibex/csr_rdata [11]),
    .Y(\i_ibex/cs_registers_i/_0592_ ),
    .B1(net559));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1747_  (.Y(\i_ibex/cs_registers_i/_0593_ ),
    .A(net559),
    .B(\i_ibex/cs_registers_i/_0228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1748_  (.A(\i_ibex/cs_registers_i/_0592_ ),
    .B_N(\i_ibex/cs_registers_i/_0593_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout963 (.X(net963),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1750_  (.S0(net496),
    .A0(\i_ibex/cs_registers_i/dcsr_q [10]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [10]),
    .A2(\i_ibex/csr_depc [10]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [10]),
    .S1(net1099),
    .X(\i_ibex/cs_registers_i/_0595_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1751_  (.Y(\i_ibex/cs_registers_i/_0596_ ),
    .A(\i_ibex/cs_registers_i/mscratch_q [10]),
    .B(net1034),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1752_  (.B(net1062),
    .C(net512),
    .A(\i_ibex/cs_registers_i/mtval_q [10]),
    .Y(\i_ibex/cs_registers_i/_0597_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1753_  (.B1(\i_ibex/cs_registers_i/_0597_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0598_ ),
    .VSS(VSS),
    .A1(net510),
    .A2(\i_ibex/cs_registers_i/_0596_ ));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1754_  (.A2(\i_ibex/cs_registers_i/_0598_ ),
    .A1(\i_ibex/cs_registers_i/_0272_ ),
    .B1(\i_ibex/cs_registers_i/_0476_ ),
    .X(\i_ibex/cs_registers_i/_0599_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1755_  (.Y(\i_ibex/cs_registers_i/_0600_ ),
    .B1(\i_ibex/cs_registers_i/_0599_ ),
    .B2(net465),
    .A2(\i_ibex/cs_registers_i/_0595_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1756_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [10]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0601_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1757_  (.Y(\i_ibex/cs_registers_i/_0602_ ),
    .B1(net1006),
    .B2(\i_ibex/cs_registers_i/_0601_ ),
    .A2(\i_ibex/cs_registers_i/_0133_ ),
    .A1(\i_ibex/csr_mtvec [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1758_  (.Y(\i_ibex/cs_registers_i/_0603_ ),
    .B1(net989),
    .B2(net23),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1759_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2026]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [42]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0604_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1760_  (.A2(net455),
    .A1(\i_ibex/csr_mepc [10]),
    .B1(\i_ibex/cs_registers_i/_0124_ ),
    .X(\i_ibex/cs_registers_i/_0605_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1761_  (.Y(\i_ibex/cs_registers_i/_0606_ ),
    .B1(\i_ibex/cs_registers_i/_0605_ ),
    .B2(\i_ibex/cs_registers_i/_0286_ ),
    .A2(\i_ibex/cs_registers_i/_0604_ ),
    .A1(net999),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1762_  (.B(\i_ibex/cs_registers_i/_0602_ ),
    .C(\i_ibex/cs_registers_i/_0603_ ),
    .A(\i_ibex/cs_registers_i/_0600_ ),
    .Y(\i_ibex/cs_registers_i/_0607_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0606_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1763_  (.A(net976),
    .B_N(\i_ibex/cs_registers_i/_0607_ ),
    .Y(\i_ibex/csr_rdata [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1764_  (.Y(\i_ibex/cs_registers_i/_0608_ ),
    .A(net691),
    .B(\i_ibex/csr_rdata [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1765_  (.Y(\i_ibex/cs_registers_i/_0609_ ),
    .A(net557),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1766_  (.B1(\i_ibex/cs_registers_i/_0609_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [10]),
    .VSS(VSS),
    .A1(net557),
    .A2(\i_ibex/cs_registers_i/_0608_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1767_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2025]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [41]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0610_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1768_  (.Y(\i_ibex/cs_registers_i/_0611_ ),
    .B1(net1002),
    .B2(\i_ibex/cs_registers_i/_0610_ ),
    .A2(net451),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1769_  (.Y(\i_ibex/cs_registers_i/_0612_ ),
    .B1(net445),
    .B2(\i_ibex/cs_registers_i/dcsr_q [9]),
    .A2(net987),
    .A1(\i_ibex/csr_mtvec [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1770_  (.A(\i_ibex/cs_registers_i/_0611_ ),
    .B(\i_ibex/cs_registers_i/_0612_ ),
    .X(\i_ibex/cs_registers_i/_0613_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1771_  (.A(\i_ibex/csr_mepc [9]),
    .B(net1066),
    .X(\i_ibex/cs_registers_i/_0614_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1772_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [9]),
    .A2(net1035),
    .Y(\i_ibex/cs_registers_i/_0615_ ),
    .B1(\i_ibex/cs_registers_i/_0614_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1773_  (.B(net1065),
    .C(net507),
    .A(\i_ibex/cs_registers_i/mtval_q [9]),
    .Y(\i_ibex/cs_registers_i/_0616_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1774_  (.B1(\i_ibex/cs_registers_i/_0616_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0617_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0615_ ));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1775_  (.A2(\i_ibex/cs_registers_i/_0617_ ),
    .A1(\i_ibex/cs_registers_i/_0272_ ),
    .B1(\i_ibex/cs_registers_i/_0476_ ),
    .X(\i_ibex/cs_registers_i/_0618_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1776_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [9]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [9]),
    .S(net1090),
    .X(\i_ibex/cs_registers_i/_0619_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1777_  (.B(\i_ibex/cs_registers_i/_0160_ ),
    .C(\i_ibex/cs_registers_i/_0619_ ),
    .A(\i_ibex/cs_registers_i/_0135_ ),
    .Y(\i_ibex/cs_registers_i/_0620_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1778_  (.A(net1098),
    .B(\i_ibex/cs_registers_i/_0058_ ),
    .Y(\i_ibex/cs_registers_i/_0621_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1779_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0622_ ),
    .A(\i_ibex/csr_depc [9]),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1780_  (.A(\i_ibex/cs_registers_i/_0622_ ),
    .B(\i_ibex/cs_registers_i/_0062_ ),
    .Y(\i_ibex/cs_registers_i/_0623_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1781_  (.A(net1095),
    .B(\i_ibex/cs_registers_i/_0056_ ),
    .C(\i_ibex/cs_registers_i/_0081_ ),
    .Y(\i_ibex/cs_registers_i/_0624_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1782_  (.B1(\i_ibex/cs_registers_i/_0624_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0625_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0621_ ),
    .A2(\i_ibex/cs_registers_i/_0623_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1783_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1993]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [9]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0626_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1784_  (.Y(\i_ibex/cs_registers_i/_0627_ ),
    .B1(net1003),
    .B2(\i_ibex/cs_registers_i/_0626_ ),
    .A2(net988),
    .A1(net24),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1785_  (.B(\i_ibex/cs_registers_i/_0625_ ),
    .C(\i_ibex/cs_registers_i/_0627_ ),
    .A(\i_ibex/cs_registers_i/_0620_ ),
    .Y(\i_ibex/cs_registers_i/_0628_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1786_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0628_ ),
    .Y(\i_ibex/cs_registers_i/_0629_ ),
    .A2(\i_ibex/cs_registers_i/_0618_ ),
    .A1(net465));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1787_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net975),
    .Y(\i_ibex/csr_rdata [9]),
    .A2(\i_ibex/cs_registers_i/_0629_ ),
    .A1(\i_ibex/cs_registers_i/_0613_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1788_  (.Y(\i_ibex/cs_registers_i/_0630_ ),
    .A(net691),
    .B(\i_ibex/csr_rdata [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1789_  (.Y(\i_ibex/cs_registers_i/_0631_ ),
    .A(net555),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1790_  (.B1(\i_ibex/cs_registers_i/_0631_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [9]),
    .VSS(VSS),
    .A1(net555),
    .A2(\i_ibex/cs_registers_i/_0630_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1791_  (.A0(\i_ibex/csr_mepc [8]),
    .A1(\i_ibex/cs_registers_i/mtval_q [8]),
    .S(net497),
    .X(\i_ibex/cs_registers_i/_0632_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1792_  (.Y(\i_ibex/cs_registers_i/_0633_ ),
    .B1(\i_ibex/cs_registers_i/_0632_ ),
    .B2(net1063),
    .A2(net1040),
    .A1(\i_ibex/cs_registers_i/mscratch_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1793_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0634_ ),
    .A(\i_ibex/cs_registers_i/_0044_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1794_  (.B1(\i_ibex/cs_registers_i/_0634_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0635_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0102_ ),
    .A2(\i_ibex/cs_registers_i/_0633_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1795_  (.B(net462),
    .C(\i_ibex/cs_registers_i/_0635_ ),
    .A(net465),
    .Y(\i_ibex/cs_registers_i/_0636_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/cs_registers_i/_1796_  (.S0(net515),
    .A0(\i_ibex/cs_registers_i/dcsr_q [8]),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [8]),
    .A2(\i_ibex/csr_depc [8]),
    .A3(\i_ibex/cs_registers_i/dscratch1_q [8]),
    .S1(net1104),
    .X(\i_ibex/cs_registers_i/_0637_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1797_  (.Y(\i_ibex/cs_registers_i/_0638_ ),
    .B1(\i_ibex/cs_registers_i/_0637_ ),
    .B2(net460),
    .A2(net987),
    .A1(\i_ibex/csr_mtvec [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1798_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1992]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [8]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0639_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1799_  (.Y(\i_ibex/cs_registers_i/_0640_ ),
    .B1(net1003),
    .B2(\i_ibex/cs_registers_i/_0639_ ),
    .A2(net988),
    .A1(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1800_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2024]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [40]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0641_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1801_  (.Y(\i_ibex/cs_registers_i/_0642_ ),
    .B1(net999),
    .B2(\i_ibex/cs_registers_i/_0641_ ),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1802_  (.B(\i_ibex/cs_registers_i/_0638_ ),
    .C(\i_ibex/cs_registers_i/_0640_ ),
    .A(\i_ibex/cs_registers_i/_0636_ ),
    .Y(\i_ibex/cs_registers_i/_0643_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0642_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1803_  (.A(net975),
    .B_N(\i_ibex/cs_registers_i/_0643_ ),
    .Y(\i_ibex/csr_rdata [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1804_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net691),
    .A2(\i_ibex/csr_rdata [8]),
    .Y(\i_ibex/cs_registers_i/_0644_ ),
    .B1(net553));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1805_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0644_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [8]),
    .A2(\i_ibex/cs_registers_i/_0228_ ),
    .A1(net553));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1806_  (.A0(\i_ibex/cs_registers_i/mscratch_q [7]),
    .A1(timer0_irq_i),
    .S(net586),
    .X(\i_ibex/cs_registers_i/_0645_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/_1807_  (.X(\i_ibex/cs_registers_i/_0646_ ),
    .A(\i_ibex/cs_registers_i/_0163_ ),
    .B(\i_ibex/cs_registers_i/mie_q [17]),
    .C(net589),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1808_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1096),
    .A2(\i_ibex/cs_registers_i/_0645_ ),
    .Y(\i_ibex/cs_registers_i/_0647_ ),
    .B1(\i_ibex/cs_registers_i/_0646_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1809_  (.A(net1093),
    .B(net588),
    .Y(\i_ibex/cs_registers_i/_0648_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1810_  (.B1(\i_ibex/cs_registers_i/_0648_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0649_ ),
    .VSS(VSS),
    .A1(net483),
    .A2(\i_ibex/cs_registers_i/mstatus_q [4]));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1811_  (.B1(\i_ibex/cs_registers_i/_0649_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0650_ ),
    .VSS(VSS),
    .A1(net483),
    .A2(\i_ibex/cs_registers_i/_0647_ ));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1812_  (.B(\i_ibex/cs_registers_i/_0071_ ),
    .C(net1031),
    .A(net465),
    .Y(\i_ibex/cs_registers_i/_0651_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0650_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1813_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2023]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [39]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0652_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1814_  (.Y(\i_ibex/cs_registers_i/_0653_ ),
    .B1(\i_ibex/cs_registers_i/_0652_ ),
    .B2(net998),
    .A2(\i_ibex/cs_registers_i/_0161_ ),
    .A1(\i_ibex/cs_registers_i/dcsr_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1815_  (.A0(\i_ibex/csr_depc [7]),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [7]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0654_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1816_  (.Y(\i_ibex/cs_registers_i/_0655_ ),
    .B1(\i_ibex/cs_registers_i/_0654_ ),
    .B2(net1062),
    .A2(\i_ibex/cs_registers_i/_0573_ ),
    .A1(\i_ibex/cs_registers_i/dscratch0_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1817_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0656_ ),
    .A(\i_ibex/cs_registers_i/_0655_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1818_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1991]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [7]),
    .S(net498),
    .X(\i_ibex/cs_registers_i/_0657_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1819_  (.Y(\i_ibex/cs_registers_i/_0658_ ),
    .B1(\i_ibex/cs_registers_i/_0657_ ),
    .B2(net1003),
    .A2(\i_ibex/cs_registers_i/_0656_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1820_  (.A0(\i_ibex/csr_mepc [7]),
    .A1(\i_ibex/cs_registers_i/mtval_q [7]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0659_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1821_  (.B(\i_ibex/cs_registers_i/_0071_ ),
    .C(\i_ibex/cs_registers_i/_0363_ ),
    .A(net473),
    .Y(\i_ibex/cs_registers_i/_0660_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0659_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1822_  (.Y(\i_ibex/cs_registers_i/_0661_ ),
    .A(\i_ibex/csr_mtvec [7]),
    .B(\i_ibex/cs_registers_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1823_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0660_ ),
    .A2(\i_ibex/cs_registers_i/_0661_ ),
    .Y(\i_ibex/cs_registers_i/_0662_ ),
    .B1(\i_ibex/cs_registers_i/_0042_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1824_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net26),
    .C1(\i_ibex/cs_registers_i/_0662_ ),
    .B1(net988),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [7]),
    .Y(\i_ibex/cs_registers_i/_0663_ ),
    .A2(net448));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1825_  (.A(\i_ibex/cs_registers_i/_0651_ ),
    .B(\i_ibex/cs_registers_i/_0653_ ),
    .C(\i_ibex/cs_registers_i/_0658_ ),
    .D(\i_ibex/cs_registers_i/_0663_ ),
    .X(\i_ibex/cs_registers_i/_0664_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1826_  (.A(net551),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0664_ ),
    .Y(\i_ibex/cs_registers_i/_0665_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/cs_registers_i/_1827_  (.A2(net633),
    .A1(net551),
    .B1(\i_ibex/cs_registers_i/_0665_ ),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout962 (.X(net962),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1829_  (.A0(\i_ibex/csr_mepc [6]),
    .A1(\i_ibex/cs_registers_i/mtval_q [6]),
    .S(net506),
    .X(\i_ibex/cs_registers_i/_0667_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1830_  (.Y(\i_ibex/cs_registers_i/_0668_ ),
    .B1(\i_ibex/cs_registers_i/_0667_ ),
    .B2(net1064),
    .A2(net1040),
    .A1(\i_ibex/cs_registers_i/mscratch_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1831_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0669_ ),
    .A(\i_ibex/cs_registers_i/_0668_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1832_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0669_ ),
    .C1(\i_ibex/cs_registers_i/_0254_ ),
    .B1(\i_ibex/cs_registers_i/_0527_ ),
    .A1(\i_ibex/csr_mtvec [6]),
    .Y(\i_ibex/cs_registers_i/_0670_ ),
    .A2(net984));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1833_  (.Y(\i_ibex/cs_registers_i/_0671_ ),
    .B1(net445),
    .B2(\i_ibex/cs_registers_i/dcsr_q [6]),
    .A2(\i_ibex/cs_registers_i/_0129_ ),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1834_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [1990]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [6]),
    .S(net500),
    .X(\i_ibex/cs_registers_i/_0672_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1835_  (.Y(\i_ibex/cs_registers_i/_0673_ ),
    .B1(net1003),
    .B2(\i_ibex/cs_registers_i/_0672_ ),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1836_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2022]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [38]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0674_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1837_  (.Y(\i_ibex/cs_registers_i/_0675_ ),
    .A(\i_ibex/csr_depc [6]),
    .B(net1064),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1838_  (.B(net1034),
    .C(net510),
    .A(\i_ibex/cs_registers_i/dscratch0_q [6]),
    .Y(\i_ibex/cs_registers_i/_0676_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1839_  (.B1(\i_ibex/cs_registers_i/_0676_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0677_ ),
    .VSS(VSS),
    .A1(net511),
    .A2(\i_ibex/cs_registers_i/_0675_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1840_  (.A(net459),
    .B(\i_ibex/cs_registers_i/_0677_ ),
    .X(\i_ibex/cs_registers_i/_0678_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1841_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0674_ ),
    .C1(\i_ibex/cs_registers_i/_0678_ ),
    .B1(net998),
    .A1(net27),
    .Y(\i_ibex/cs_registers_i/_0679_ ),
    .A2(net988));
 sg13g2_and4_2 \i_ibex/cs_registers_i/_1842_  (.A(\i_ibex/cs_registers_i/_0670_ ),
    .B(\i_ibex/cs_registers_i/_0671_ ),
    .C(\i_ibex/cs_registers_i/_0673_ ),
    .D(\i_ibex/cs_registers_i/_0679_ ),
    .X(\i_ibex/cs_registers_i/_0680_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_1843_  (.A(\i_ibex/alu_operand_a_ex [6]),
    .B(\i_ibex/cs_registers_i/_0153_ ),
    .C(\i_ibex/cs_registers_i/_0680_ ),
    .Y(\i_ibex/cs_registers_i/_0681_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1844_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/cs_registers_i/_0681_ ),
    .Y(\i_ibex/cs_registers_i/_0682_ ),
    .A2(net634),
    .A1(\i_ibex/alu_operand_a_ex [6]));
 sg13g2_inv_4 \i_ibex/cs_registers_i/_1845_  (.A(\i_ibex/cs_registers_i/_0682_ ),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1846_  (.Y(\i_ibex/cs_registers_i/_0683_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [28]),
    .A2(net990),
    .A1(net28),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1847_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2044]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [60]),
    .S(net505),
    .X(\i_ibex/cs_registers_i/_0684_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1848_  (.A(net1103),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [28]),
    .Y(\i_ibex/cs_registers_i/_0685_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1849_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [28]),
    .A2(net1103),
    .Y(\i_ibex/cs_registers_i/_0686_ ),
    .B1(\i_ibex/cs_registers_i/_0685_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1850_  (.B(net1036),
    .C(net512),
    .A(\i_ibex/cs_registers_i/dscratch0_q [28]),
    .Y(\i_ibex/cs_registers_i/_0687_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1851_  (.B1(\i_ibex/cs_registers_i/_0687_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0688_ ),
    .VSS(VSS),
    .A1(net510),
    .A2(\i_ibex/cs_registers_i/_0686_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1852_  (.Y(\i_ibex/cs_registers_i/_0689_ ),
    .B1(\i_ibex/cs_registers_i/_0688_ ),
    .B2(net460),
    .A2(\i_ibex/cs_registers_i/_0684_ ),
    .A1(net1000),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1853_  (.A(\i_ibex/cs_registers_i/_0683_ ),
    .B(\i_ibex/cs_registers_i/_0689_ ),
    .X(\i_ibex/cs_registers_i/_0690_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1854_  (.A0(\i_ibex/csr_mepc [28]),
    .A1(\i_ibex/cs_registers_i/mtval_q [28]),
    .S(net499),
    .X(\i_ibex/cs_registers_i/_0691_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1855_  (.Y(\i_ibex/cs_registers_i/_0692_ ),
    .B1(\i_ibex/cs_registers_i/_0691_ ),
    .B2(net1070),
    .A2(\i_ibex/cs_registers_i/_0026_ ),
    .A1(\i_ibex/cs_registers_i/mscratch_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1856_  (.Y(\i_ibex/cs_registers_i/_0693_ ),
    .A(irqs_i[12]),
    .B(net457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1857_  (.B1(\i_ibex/cs_registers_i/_0693_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0694_ ),
    .VSS(VSS),
    .A1(net1033),
    .A2(\i_ibex/cs_registers_i/_0692_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1858_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [28]),
    .C1(net982),
    .B1(net446),
    .A1(\i_ibex/cs_registers_i/mie_q [12]),
    .Y(\i_ibex/cs_registers_i/_0695_ ),
    .A2(net436));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_1859_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2012]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [28]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0696_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1860_  (.Y(\i_ibex/cs_registers_i/_0697_ ),
    .B1(net1004),
    .B2(\i_ibex/cs_registers_i/_0696_ ),
    .A2(net985),
    .A1(\i_ibex/csr_mtvec [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1861_  (.Y(\i_ibex/cs_registers_i/_0698_ ),
    .A(\i_ibex/cs_registers_i/_0695_ ),
    .B(\i_ibex/cs_registers_i/_0697_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1862_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net454),
    .A2(\i_ibex/cs_registers_i/_0694_ ),
    .Y(\i_ibex/cs_registers_i/_0699_ ),
    .B1(\i_ibex/cs_registers_i/_0698_ ));
 sg13g2_a21oi_2 \i_ibex/cs_registers_i/_1863_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net977),
    .Y(\i_ibex/csr_rdata [28]),
    .A2(\i_ibex/cs_registers_i/_0699_ ),
    .A1(\i_ibex/cs_registers_i/_0690_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1864_  (.Y(\i_ibex/cs_registers_i/_0700_ ),
    .A(net691),
    .B(\i_ibex/csr_rdata [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1865_  (.Y(\i_ibex/cs_registers_i/_0701_ ),
    .A(net539),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1866_  (.B1(\i_ibex/cs_registers_i/_0701_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [28]),
    .VSS(VSS),
    .A1(net539),
    .A2(\i_ibex/cs_registers_i/_0700_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_1867_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0702_ ),
    .B(\i_ibex/cs_registers_i/_0016_ ),
    .A(net1032));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1868_  (.Y(\i_ibex/cs_registers_i/_0703_ ),
    .B1(net453),
    .B2(\i_ibex/cs_registers_i/mtval_q [27]),
    .A2(\i_ibex/cs_registers_i/_0127_ ),
    .A1(\i_ibex/cs_registers_i/dscratch1_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_1869_  (.A(\i_ibex/cs_registers_i/_0702_ ),
    .B(\i_ibex/cs_registers_i/_0703_ ),
    .Y(\i_ibex/cs_registers_i/_0704_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1870_  (.A(\i_ibex/cs_registers_i/mie_q [11]),
    .B(net436),
    .X(\i_ibex/cs_registers_i/_0705_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1871_  (.A0(\i_ibex/cs_registers_i/mscratch_q [27]),
    .A1(irqs_i[11]),
    .S(net586),
    .X(\i_ibex/cs_registers_i/_0706_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1872_  (.Y(\i_ibex/cs_registers_i/_0707_ ),
    .B1(\i_ibex/cs_registers_i/_0706_ ),
    .B2(net1039),
    .A2(\i_ibex/cs_registers_i/_0362_ ),
    .A1(\i_ibex/csr_mepc [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1873_  (.A(\i_ibex/cs_registers_i/_0707_ ),
    .B_N(\i_ibex/cs_registers_i/_0566_ ),
    .Y(\i_ibex/cs_registers_i/_0708_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1874_  (.Y(\i_ibex/cs_registers_i/_0709_ ),
    .B1(\i_ibex/cs_registers_i/_0135_ ),
    .B2(\i_ibex/cs_registers_i/dscratch0_q [27]),
    .A2(\i_ibex/cs_registers_i/_0286_ ),
    .A1(\i_ibex/csr_depc [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1875_  (.A(\i_ibex/cs_registers_i/_0709_ ),
    .B_N(\i_ibex/cs_registers_i/_0127_ ),
    .Y(\i_ibex/cs_registers_i/_0710_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/cs_registers_i/_1876_  (.A(\i_ibex/cs_registers_i/_0254_ ),
    .B(\i_ibex/cs_registers_i/_0705_ ),
    .C(\i_ibex/cs_registers_i/_0708_ ),
    .D(\i_ibex/cs_registers_i/_0710_ ),
    .X(\i_ibex/cs_registers_i/_0711_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1877_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2011]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [27]),
    .S(net502),
    .X(\i_ibex/cs_registers_i/_0712_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1878_  (.Y(\i_ibex/cs_registers_i/_0713_ ),
    .B1(\i_ibex/cs_registers_i/_0712_ ),
    .B2(net1006),
    .A2(net445),
    .A1(\i_ibex/cs_registers_i/dcsr_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_1879_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0714_ ),
    .A(\i_ibex/cs_registers_i/_0713_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1880_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2043]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [59]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0715_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1881_  (.Y(\i_ibex/cs_registers_i/_0716_ ),
    .B1(net1001),
    .B2(\i_ibex/cs_registers_i/_0715_ ),
    .A2(net987),
    .A1(\i_ibex/csr_mtvec [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1882_  (.Y(\i_ibex/cs_registers_i/_0717_ ),
    .B1(net991),
    .B2(net29),
    .A2(net448),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1883_  (.Y(\i_ibex/cs_registers_i/_0718_ ),
    .A(\i_ibex/cs_registers_i/_0716_ ),
    .B(\i_ibex/cs_registers_i/_0717_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_1884_  (.A(\i_ibex/cs_registers_i/_0704_ ),
    .B(\i_ibex/cs_registers_i/_0711_ ),
    .C(\i_ibex/cs_registers_i/_0714_ ),
    .Y(\i_ibex/cs_registers_i/_0719_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0718_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_1885_  (.A(net534),
    .B(\i_ibex/cs_registers_i/_0295_ ),
    .C(net979),
    .D(\i_ibex/cs_registers_i/_0719_ ),
    .Y(\i_ibex/cs_registers_i/_0720_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_1886_  (.A2(net633),
    .A1(net534),
    .B1(\i_ibex/cs_registers_i/_0720_ ),
    .X(\i_ibex/cs_registers_i/csr_wdata_int [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(net962),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1888_  (.A(\i_ibex/csr_mepc [26]),
    .B(net1069),
    .X(\i_ibex/cs_registers_i/_0722_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1889_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [26]),
    .A2(net1037),
    .Y(\i_ibex/cs_registers_i/_0723_ ),
    .B1(\i_ibex/cs_registers_i/_0722_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1890_  (.B(net1070),
    .C(net514),
    .A(\i_ibex/cs_registers_i/mtval_q [26]),
    .Y(\i_ibex/cs_registers_i/_0724_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1891_  (.B1(\i_ibex/cs_registers_i/_0724_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0725_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0723_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1892_  (.Y(\i_ibex/cs_registers_i/_0726_ ),
    .B1(\i_ibex/cs_registers_i/_0725_ ),
    .B2(net1042),
    .A2(net456),
    .A1(irqs_i[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1893_  (.Y(\i_ibex/cs_registers_i/_0727_ ),
    .B(net454),
    .A_N(\i_ibex/cs_registers_i/_0726_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1894_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/csr_mtvec [26]),
    .C1(net982),
    .B1(net985),
    .A1(\i_ibex/cs_registers_i/mie_q [10]),
    .Y(\i_ibex/cs_registers_i/_0728_ ),
    .A2(net437));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1895_  (.Y(\i_ibex/cs_registers_i/_0729_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [26]),
    .A2(net990),
    .A1(net30),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1896_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2042]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [58]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0730_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1897_  (.Y(\i_ibex/cs_registers_i/_0731_ ),
    .B1(net1000),
    .B2(\i_ibex/cs_registers_i/_0730_ ),
    .A2(net447),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1898_  (.A(net1102),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [26]),
    .Y(\i_ibex/cs_registers_i/_0732_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1899_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [26]),
    .A2(net1101),
    .Y(\i_ibex/cs_registers_i/_0733_ ),
    .B1(\i_ibex/cs_registers_i/_0732_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1900_  (.B(net1036),
    .C(net509),
    .A(\i_ibex/cs_registers_i/dscratch0_q [26]),
    .Y(\i_ibex/cs_registers_i/_0734_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1901_  (.B1(\i_ibex/cs_registers_i/_0734_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0735_ ),
    .VSS(VSS),
    .A1(net514),
    .A2(\i_ibex/cs_registers_i/_0733_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1902_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [26]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0736_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1903_  (.Y(\i_ibex/cs_registers_i/_0737_ ),
    .B1(\i_ibex/cs_registers_i/_0736_ ),
    .B2(net1004),
    .A2(\i_ibex/cs_registers_i/_0735_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1904_  (.A(\i_ibex/cs_registers_i/_0731_ ),
    .B(\i_ibex/cs_registers_i/_0737_ ),
    .X(\i_ibex/cs_registers_i/_0738_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1905_  (.B(\i_ibex/cs_registers_i/_0728_ ),
    .C(\i_ibex/cs_registers_i/_0729_ ),
    .A(\i_ibex/cs_registers_i/_0727_ ),
    .Y(\i_ibex/cs_registers_i/_0739_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0738_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1906_  (.A(net978),
    .B_N(\i_ibex/cs_registers_i/_0739_ ),
    .Y(\i_ibex/csr_rdata [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1907_  (.Y(\i_ibex/cs_registers_i/_0740_ ),
    .A(net691),
    .B(\i_ibex/csr_rdata [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1908_  (.Y(\i_ibex/cs_registers_i/_0741_ ),
    .A(\i_ibex/alu_operand_a_ex [26]),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1909_  (.B1(\i_ibex/cs_registers_i/_0741_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [26]),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_a_ex [26]),
    .A2(\i_ibex/cs_registers_i/_0740_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1910_  (.A(\i_ibex/csr_mepc [25]),
    .B(net1069),
    .X(\i_ibex/cs_registers_i/_0742_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1911_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [25]),
    .A2(net1037),
    .Y(\i_ibex/cs_registers_i/_0743_ ),
    .B1(\i_ibex/cs_registers_i/_0742_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1912_  (.B(net1070),
    .C(net514),
    .A(\i_ibex/cs_registers_i/mtval_q [25]),
    .Y(\i_ibex/cs_registers_i/_0744_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1913_  (.B1(\i_ibex/cs_registers_i/_0744_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0745_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0743_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1914_  (.Y(\i_ibex/cs_registers_i/_0746_ ),
    .B1(\i_ibex/cs_registers_i/_0745_ ),
    .B2(net1042),
    .A2(net456),
    .A1(irqs_i[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1915_  (.Y(\i_ibex/cs_registers_i/_0747_ ),
    .B(net454),
    .A_N(\i_ibex/cs_registers_i/_0746_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1916_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/csr_mtvec [25]),
    .C1(net982),
    .B1(net985),
    .A1(\i_ibex/cs_registers_i/mie_q [9]),
    .Y(\i_ibex/cs_registers_i/_0748_ ),
    .A2(net437));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1917_  (.Y(\i_ibex/cs_registers_i/_0749_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [25]),
    .A2(net990),
    .A1(net31),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1918_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2041]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [57]),
    .S(net504),
    .X(\i_ibex/cs_registers_i/_0750_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1919_  (.Y(\i_ibex/cs_registers_i/_0751_ ),
    .B1(net1000),
    .B2(\i_ibex/cs_registers_i/_0750_ ),
    .A2(net447),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1920_  (.A(net1103),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [25]),
    .Y(\i_ibex/cs_registers_i/_0752_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1921_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [25]),
    .A2(net1104),
    .Y(\i_ibex/cs_registers_i/_0753_ ),
    .B1(\i_ibex/cs_registers_i/_0752_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1922_  (.B(net1036),
    .C(net509),
    .A(\i_ibex/cs_registers_i/dscratch0_q [25]),
    .Y(\i_ibex/cs_registers_i/_0754_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1923_  (.B1(\i_ibex/cs_registers_i/_0754_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0755_ ),
    .VSS(VSS),
    .A1(net514),
    .A2(\i_ibex/cs_registers_i/_0753_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1924_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [25]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0756_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1925_  (.Y(\i_ibex/cs_registers_i/_0757_ ),
    .B1(\i_ibex/cs_registers_i/_0756_ ),
    .B2(net1004),
    .A2(\i_ibex/cs_registers_i/_0755_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1926_  (.A(\i_ibex/cs_registers_i/_0751_ ),
    .B(\i_ibex/cs_registers_i/_0757_ ),
    .X(\i_ibex/cs_registers_i/_0758_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1927_  (.B(\i_ibex/cs_registers_i/_0748_ ),
    .C(\i_ibex/cs_registers_i/_0749_ ),
    .A(\i_ibex/cs_registers_i/_0747_ ),
    .Y(\i_ibex/cs_registers_i/_0759_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0758_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1928_  (.A(net977),
    .B_N(\i_ibex/cs_registers_i/_0759_ ),
    .Y(\i_ibex/csr_rdata [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1929_  (.Y(\i_ibex/cs_registers_i/_0760_ ),
    .A(net690),
    .B(\i_ibex/csr_rdata [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1930_  (.Y(\i_ibex/cs_registers_i/_0761_ ),
    .A(net530),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1931_  (.B1(\i_ibex/cs_registers_i/_0761_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [25]),
    .VSS(VSS),
    .A1(net530),
    .A2(\i_ibex/cs_registers_i/_0760_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1932_  (.A(\i_ibex/csr_mepc [24]),
    .B(net1069),
    .X(\i_ibex/cs_registers_i/_0762_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1933_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [24]),
    .A2(net1039),
    .Y(\i_ibex/cs_registers_i/_0763_ ),
    .B1(\i_ibex/cs_registers_i/_0762_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1934_  (.B(net1069),
    .C(net514),
    .A(\i_ibex/cs_registers_i/mtval_q [24]),
    .Y(\i_ibex/cs_registers_i/_0764_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1935_  (.B1(\i_ibex/cs_registers_i/_0764_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0765_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0763_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1936_  (.Y(\i_ibex/cs_registers_i/_0766_ ),
    .B1(\i_ibex/cs_registers_i/_0765_ ),
    .B2(net1042),
    .A2(net456),
    .A1(irqs_i[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1937_  (.Y(\i_ibex/cs_registers_i/_0767_ ),
    .B(net453),
    .A_N(\i_ibex/cs_registers_i/_0766_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1938_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/csr_mtvec [24]),
    .C1(net982),
    .B1(net985),
    .A1(\i_ibex/cs_registers_i/mie_q [8]),
    .Y(\i_ibex/cs_registers_i/_0768_ ),
    .A2(net436));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1939_  (.Y(\i_ibex/cs_registers_i/_0769_ ),
    .B1(net451),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [24]),
    .A2(net990),
    .A1(net32),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1940_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2040]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [56]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0770_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1941_  (.Y(\i_ibex/cs_registers_i/_0771_ ),
    .B1(net1000),
    .B2(\i_ibex/cs_registers_i/_0770_ ),
    .A2(net447),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1942_  (.A(net1102),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [24]),
    .Y(\i_ibex/cs_registers_i/_0772_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1943_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [24]),
    .A2(net1102),
    .Y(\i_ibex/cs_registers_i/_0773_ ),
    .B1(\i_ibex/cs_registers_i/_0772_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1944_  (.B(net1036),
    .C(net509),
    .A(\i_ibex/cs_registers_i/dscratch0_q [24]),
    .Y(\i_ibex/cs_registers_i/_0774_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1945_  (.B1(\i_ibex/cs_registers_i/_0774_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0775_ ),
    .VSS(VSS),
    .A1(net514),
    .A2(\i_ibex/cs_registers_i/_0773_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1946_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [24]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0776_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1947_  (.Y(\i_ibex/cs_registers_i/_0777_ ),
    .B1(\i_ibex/cs_registers_i/_0776_ ),
    .B2(net1004),
    .A2(\i_ibex/cs_registers_i/_0775_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1948_  (.A(\i_ibex/cs_registers_i/_0771_ ),
    .B(\i_ibex/cs_registers_i/_0777_ ),
    .X(\i_ibex/cs_registers_i/_0778_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1949_  (.B(\i_ibex/cs_registers_i/_0768_ ),
    .C(\i_ibex/cs_registers_i/_0769_ ),
    .A(\i_ibex/cs_registers_i/_0767_ ),
    .Y(\i_ibex/cs_registers_i/_0779_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0778_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1950_  (.A(net977),
    .B_N(\i_ibex/cs_registers_i/_0779_ ),
    .Y(\i_ibex/csr_rdata [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1951_  (.Y(\i_ibex/cs_registers_i/_0780_ ),
    .A(net690),
    .B(\i_ibex/csr_rdata [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1952_  (.Y(\i_ibex/cs_registers_i/_0781_ ),
    .A(net528),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1953_  (.B1(\i_ibex/cs_registers_i/_0781_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [24]),
    .VSS(VSS),
    .A1(net528),
    .A2(\i_ibex/cs_registers_i/_0780_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1954_  (.A(\i_ibex/csr_mepc [23]),
    .B(net1069),
    .X(\i_ibex/cs_registers_i/_0782_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1955_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [23]),
    .A2(net1037),
    .Y(\i_ibex/cs_registers_i/_0783_ ),
    .B1(\i_ibex/cs_registers_i/_0782_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1956_  (.B(net1070),
    .C(net514),
    .A(\i_ibex/cs_registers_i/mtval_q [23]),
    .Y(\i_ibex/cs_registers_i/_0784_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1957_  (.B1(\i_ibex/cs_registers_i/_0784_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0785_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0783_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1958_  (.Y(\i_ibex/cs_registers_i/_0786_ ),
    .B1(\i_ibex/cs_registers_i/_0785_ ),
    .B2(net1042),
    .A2(net456),
    .A1(irqs_i[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1959_  (.Y(\i_ibex/cs_registers_i/_0787_ ),
    .B(net453),
    .A_N(\i_ibex/cs_registers_i/_0786_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1960_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/csr_mtvec [23]),
    .C1(net982),
    .B1(net985),
    .A1(\i_ibex/cs_registers_i/mie_q [7]),
    .Y(\i_ibex/cs_registers_i/_0788_ ),
    .A2(net436));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1961_  (.Y(\i_ibex/cs_registers_i/_0789_ ),
    .B1(net450),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [23]),
    .A2(\i_ibex/cs_registers_i/_0125_ ),
    .A1(net33),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1962_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2039]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [55]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0790_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1963_  (.Y(\i_ibex/cs_registers_i/_0791_ ),
    .B1(net1000),
    .B2(\i_ibex/cs_registers_i/_0790_ ),
    .A2(net447),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1964_  (.A(net1103),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [23]),
    .Y(\i_ibex/cs_registers_i/_0792_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1965_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [23]),
    .A2(net1102),
    .Y(\i_ibex/cs_registers_i/_0793_ ),
    .B1(\i_ibex/cs_registers_i/_0792_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1966_  (.B(net1036),
    .C(net509),
    .A(\i_ibex/cs_registers_i/dscratch0_q [23]),
    .Y(\i_ibex/cs_registers_i/_0794_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1967_  (.B1(\i_ibex/cs_registers_i/_0794_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0795_ ),
    .VSS(VSS),
    .A1(net514),
    .A2(\i_ibex/cs_registers_i/_0793_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1968_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2007]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [23]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0796_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1969_  (.Y(\i_ibex/cs_registers_i/_0797_ ),
    .B1(\i_ibex/cs_registers_i/_0796_ ),
    .B2(net1004),
    .A2(\i_ibex/cs_registers_i/_0795_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1970_  (.A(\i_ibex/cs_registers_i/_0791_ ),
    .B(\i_ibex/cs_registers_i/_0797_ ),
    .X(\i_ibex/cs_registers_i/_0798_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1971_  (.B(\i_ibex/cs_registers_i/_0788_ ),
    .C(\i_ibex/cs_registers_i/_0789_ ),
    .A(\i_ibex/cs_registers_i/_0787_ ),
    .Y(\i_ibex/cs_registers_i/_0799_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0798_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1972_  (.A(net977),
    .B_N(\i_ibex/cs_registers_i/_0799_ ),
    .Y(\i_ibex/csr_rdata [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1973_  (.Y(\i_ibex/cs_registers_i/_0800_ ),
    .A(net689),
    .B(\i_ibex/csr_rdata [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1974_  (.Y(\i_ibex/cs_registers_i/_0801_ ),
    .A(net594),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1975_  (.B1(\i_ibex/cs_registers_i/_0801_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [23]),
    .VSS(VSS),
    .A1(net594),
    .A2(\i_ibex/cs_registers_i/_0800_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1976_  (.A(\i_ibex/csr_mepc [22]),
    .B(net1069),
    .X(\i_ibex/cs_registers_i/_0802_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1977_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mscratch_q [22]),
    .A2(net1037),
    .Y(\i_ibex/cs_registers_i/_0803_ ),
    .B1(\i_ibex/cs_registers_i/_0802_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1978_  (.B(net1070),
    .C(net513),
    .A(\i_ibex/cs_registers_i/mtval_q [22]),
    .Y(\i_ibex/cs_registers_i/_0804_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1979_  (.B1(\i_ibex/cs_registers_i/_0804_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0805_ ),
    .VSS(VSS),
    .A1(net513),
    .A2(\i_ibex/cs_registers_i/_0803_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1980_  (.Y(\i_ibex/cs_registers_i/_0806_ ),
    .B1(\i_ibex/cs_registers_i/_0805_ ),
    .B2(net1042),
    .A2(net456),
    .A1(irqs_i[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_1981_  (.Y(\i_ibex/cs_registers_i/_0807_ ),
    .B(net453),
    .A_N(\i_ibex/cs_registers_i/_0806_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_1982_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/csr_mtvec [22]),
    .C1(net982),
    .B1(net985),
    .A1(\i_ibex/cs_registers_i/mie_q [6]),
    .Y(\i_ibex/cs_registers_i/_0808_ ),
    .A2(net436));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1983_  (.Y(\i_ibex/cs_registers_i/_0809_ ),
    .B1(net450),
    .B2(\i_ibex/cs_registers_i/dscratch1_q [22]),
    .A2(net991),
    .A1(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1984_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2038]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [54]),
    .S(net503),
    .X(\i_ibex/cs_registers_i/_0810_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1985_  (.Y(\i_ibex/cs_registers_i/_0811_ ),
    .B1(net1000),
    .B2(\i_ibex/cs_registers_i/_0810_ ),
    .A2(net447),
    .A1(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_1986_  (.A(net1103),
    .B_N(\i_ibex/cs_registers_i/dcsr_q [22]),
    .Y(\i_ibex/cs_registers_i/_0812_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_1987_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_depc [22]),
    .A2(net1102),
    .Y(\i_ibex/cs_registers_i/_0813_ ),
    .B1(\i_ibex/cs_registers_i/_0812_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_1988_  (.B(net1037),
    .C(net509),
    .A(\i_ibex/cs_registers_i/dscratch0_q [22]),
    .Y(\i_ibex/cs_registers_i/_0814_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1989_  (.B1(\i_ibex/cs_registers_i/_0814_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0815_ ),
    .VSS(VSS),
    .A1(net508),
    .A2(\i_ibex/cs_registers_i/_0813_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_1990_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2006]),
    .A1(\i_ibex/cs_registers_i/minstret_raw [22]),
    .S(net501),
    .X(\i_ibex/cs_registers_i/_0816_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_1991_  (.Y(\i_ibex/cs_registers_i/_0817_ ),
    .B1(\i_ibex/cs_registers_i/_0816_ ),
    .B2(net1004),
    .A2(\i_ibex/cs_registers_i/_0815_ ),
    .A1(net458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_1992_  (.A(\i_ibex/cs_registers_i/_0811_ ),
    .B(\i_ibex/cs_registers_i/_0817_ ),
    .X(\i_ibex/cs_registers_i/_0818_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_1993_  (.B(\i_ibex/cs_registers_i/_0808_ ),
    .C(\i_ibex/cs_registers_i/_0809_ ),
    .A(\i_ibex/cs_registers_i/_0807_ ),
    .Y(\i_ibex/cs_registers_i/_0819_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0818_ ));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_1994_  (.A(net977),
    .B_N(\i_ibex/cs_registers_i/_0819_ ),
    .Y(\i_ibex/csr_rdata [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1995_  (.Y(\i_ibex/cs_registers_i/_0820_ ),
    .A(net689),
    .B(\i_ibex/csr_rdata [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_1996_  (.Y(\i_ibex/cs_registers_i/_0821_ ),
    .A(\i_ibex/alu_operand_a_ex [22]),
    .B(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_1997_  (.B1(\i_ibex/cs_registers_i/_0821_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/csr_wdata_int [22]),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_a_ex [22]),
    .A2(\i_ibex/cs_registers_i/_0820_ ));
 sg13g2_buf_2 fanout960 (.A(\i_ibex/cs_registers_i/csr_wdata_int [15]),
    .X(net960),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_1999_  (.A(net979),
    .B(\i_ibex/cs_registers_i/_0354_ ),
    .Y(\i_ibex/csr_rdata [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2000_  (.A(net979),
    .B(\i_ibex/cs_registers_i/_0389_ ),
    .Y(\i_ibex/csr_rdata [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2001_  (.A(net979),
    .B(\i_ibex/cs_registers_i/_0487_ ),
    .Y(\i_ibex/csr_rdata [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2002_  (.A(net980),
    .B(\i_ibex/cs_registers_i/_0504_ ),
    .Y(\i_ibex/csr_rdata [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2003_  (.A(net979),
    .B(\i_ibex/cs_registers_i/_0522_ ),
    .Y(\i_ibex/csr_rdata [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2004_  (.VDD(VDD),
    .Y(\i_ibex/csr_rdata [12]),
    .A(\i_ibex/cs_registers_i/_0546_ ),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2005_  (.A(net980),
    .B(\i_ibex/cs_registers_i/_0664_ ),
    .Y(\i_ibex/csr_rdata [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2006_  (.A(net976),
    .B(\i_ibex/cs_registers_i/_0680_ ),
    .Y(\i_ibex/csr_rdata [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2007_  (.A(net976),
    .B(\i_ibex/cs_registers_i/_0193_ ),
    .Y(\i_ibex/csr_rdata [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2008_  (.A(net976),
    .B(\i_ibex/cs_registers_i/_0311_ ),
    .Y(\i_ibex/csr_rdata [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2009_  (.A(net976),
    .B(\i_ibex/cs_registers_i/_0334_ ),
    .Y(\i_ibex/csr_rdata [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/_2010_  (.A(net979),
    .B(\i_ibex/cs_registers_i/_0719_ ),
    .Y(\i_ibex/csr_rdata [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2011_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0287_ ),
    .A2(net1032),
    .Y(\i_ibex/cs_registers_i/_0823_ ),
    .B1(\i_ibex/cs_registers_i/_0032_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2012_  (.B(\i_ibex/cs_registers_i/_0120_ ),
    .C(\i_ibex/cs_registers_i/_0823_ ),
    .A(net464),
    .Y(\i_ibex/cs_registers_i/_0824_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_2013_  (.A(net786),
    .B_N(\i_ibex/csr_addr [8]),
    .Y(\i_ibex/cs_registers_i/_0825_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2014_  (.Y(\i_ibex/cs_registers_i/_0826_ ),
    .A(\i_ibex/csr_addr [9]),
    .B(\i_ibex/cs_registers_i/_0825_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2015_  (.Y(\i_ibex/cs_registers_i/_0827_ ),
    .A(net785),
    .B(\i_ibex/cs_registers_i/_0826_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2016_  (.B1(\i_ibex/cs_registers_i/_0827_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0828_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_addr [9]),
    .A2(\i_ibex/cs_registers_i/_0825_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_2017_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0829_ ),
    .B(\i_ibex/csr_op [0]),
    .A(net689));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2018_  (.B(\i_ibex/csr_addr [11]),
    .C(\i_ibex/cs_registers_i/_0829_ ),
    .A(\i_ibex/csr_addr [10]),
    .Y(\i_ibex/cs_registers_i/_0830_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2019_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0831_ ),
    .A(net784),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2020_  (.Y(\i_ibex/cs_registers_i/_0832_ ),
    .A(\i_ibex/cs_registers_i/_0831_ ),
    .B(net459),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2021_  (.B(\i_ibex/cs_registers_i/_0828_ ),
    .C(\i_ibex/cs_registers_i/_0830_ ),
    .A(\i_ibex/cs_registers_i/_0824_ ),
    .Y(\i_ibex/cs_registers_i/_0833_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0832_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2022_  (.A(net506),
    .B(net588),
    .X(\i_ibex/cs_registers_i/_0834_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2023_  (.Y(\i_ibex/cs_registers_i/_0835_ ),
    .A(net1089),
    .B(\i_ibex/cs_registers_i/_0834_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2024_  (.A(net483),
    .B(net1092),
    .X(\i_ibex/cs_registers_i/_0836_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2025_  (.A(net483),
    .B(net1067),
    .C(\i_ibex/cs_registers_i/_0010_ ),
    .Y(\i_ibex/cs_registers_i/_0837_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2026_  (.Y(\i_ibex/cs_registers_i/_0838_ ),
    .B1(\i_ibex/cs_registers_i/_0837_ ),
    .B2(\i_ibex/cs_registers_i/_0834_ ),
    .A2(\i_ibex/cs_registers_i/_0836_ ),
    .A1(\i_ibex/cs_registers_i/_0835_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2027_  (.B(\i_ibex/cs_registers_i/_0621_ ),
    .C(\i_ibex/cs_registers_i/_0057_ ),
    .A(net1099),
    .Y(\i_ibex/cs_registers_i/_0839_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0053_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2028_  (.B1(\i_ibex/cs_registers_i/_0839_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0840_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0038_ ),
    .A2(\i_ibex/cs_registers_i/_0838_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2029_  (.B1(\i_ibex/cs_registers_i/_0032_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0841_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0324_ ),
    .A2(\i_ibex/cs_registers_i/_0834_ ));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_2030_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0324_ ),
    .C1(\i_ibex/cs_registers_i/_0841_ ),
    .B1(\i_ibex/cs_registers_i/_0834_ ),
    .A1(\i_ibex/cs_registers_i/_0287_ ),
    .Y(\i_ibex/cs_registers_i/_0842_ ),
    .A2(\i_ibex/cs_registers_i/_0017_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2031_  (.Y(\i_ibex/cs_registers_i/_0843_ ),
    .A(\i_ibex/cs_registers_i/_0120_ ),
    .B(\i_ibex/cs_registers_i/_0107_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_2032_  (.A(net1088),
    .B(\i_ibex/cs_registers_i/_0047_ ),
    .C(\i_ibex/cs_registers_i/_0102_ ),
    .D(\i_ibex/cs_registers_i/_0103_ ),
    .Y(\i_ibex/cs_registers_i/_0844_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_2033_  (.A(net1097),
    .B(\i_ibex/cs_registers_i/_0324_ ),
    .C(\i_ibex/cs_registers_i/_0066_ ),
    .D(\i_ibex/cs_registers_i/_0134_ ),
    .Y(\i_ibex/cs_registers_i/_0845_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2034_  (.B1(\i_ibex/cs_registers_i/_0013_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0846_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0844_ ),
    .A2(\i_ibex/cs_registers_i/_0845_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2035_  (.B1(\i_ibex/cs_registers_i/_0846_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0847_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0842_ ),
    .A2(\i_ibex/cs_registers_i/_0843_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2036_  (.A0(net1067),
    .A1(\i_ibex/cs_registers_i/_0016_ ),
    .S(\i_ibex/cs_registers_i/_0324_ ),
    .X(\i_ibex/cs_registers_i/_0848_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2037_  (.A(net586),
    .B(\i_ibex/cs_registers_i/_0329_ ),
    .C(\i_ibex/cs_registers_i/_0848_ ),
    .Y(\i_ibex/cs_registers_i/_0849_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2038_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1093),
    .A2(net588),
    .Y(\i_ibex/cs_registers_i/_0850_ ),
    .B1(net1091));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_2039_  (.A(net483),
    .B(net1065),
    .C(net518),
    .D(net1088),
    .Y(\i_ibex/cs_registers_i/_0851_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2040_  (.B1(\i_ibex/cs_registers_i/_0851_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0852_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0648_ ),
    .A2(\i_ibex/cs_registers_i/_0850_ ));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2041_  (.A(net1097),
    .B(\i_ibex/cs_registers_i/_0042_ ),
    .C(\i_ibex/cs_registers_i/_0852_ ),
    .Y(\i_ibex/cs_registers_i/_0853_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2042_  (.Y(\i_ibex/cs_registers_i/_0854_ ),
    .A(net1106),
    .B(net1091),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/_2043_  (.A(net1041),
    .B(\i_ibex/cs_registers_i/_0040_ ),
    .C(\i_ibex/cs_registers_i/_0554_ ),
    .D(\i_ibex/cs_registers_i/_0854_ ),
    .X(\i_ibex/cs_registers_i/_0855_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2044_  (.Y(\i_ibex/cs_registers_i/_0856_ ),
    .B(\i_ibex/cs_registers_i/_0287_ ),
    .A_N(\i_ibex/cs_registers_i/_0061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_2045_  (.A(\i_ibex/csr_addr [11]),
    .B_N(net1098),
    .Y(\i_ibex/cs_registers_i/_0857_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2046_  (.B(\i_ibex/cs_registers_i/_0052_ ),
    .C(net473),
    .A(net1042),
    .Y(\i_ibex/cs_registers_i/_0858_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0857_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2047_  (.B1(net619),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0859_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0856_ ),
    .A2(\i_ibex/cs_registers_i/_0858_ ));
 sg13g2_or4_1 \i_ibex/cs_registers_i/_2048_  (.A(\i_ibex/cs_registers_i/_0849_ ),
    .B(\i_ibex/cs_registers_i/_0853_ ),
    .C(\i_ibex/cs_registers_i/_0855_ ),
    .D(\i_ibex/cs_registers_i/_0859_ ),
    .X(\i_ibex/cs_registers_i/_0860_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_2049_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net464),
    .C1(\i_ibex/cs_registers_i/_0860_ ),
    .B1(\i_ibex/cs_registers_i/_0847_ ),
    .A1(\i_ibex/cs_registers_i/_0163_ ),
    .Y(\i_ibex/cs_registers_i/_0861_ ),
    .A2(\i_ibex/cs_registers_i/_0840_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2050_  (.A(\i_ibex/cs_registers_i/_0051_ ),
    .B(\i_ibex/cs_registers_i/_0077_ ),
    .Y(\i_ibex/cs_registers_i/_0862_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2051_  (.Y(\i_ibex/cs_registers_i/_0863_ ),
    .A(\i_ibex/csr_op_en ),
    .B(\i_ibex/cs_registers_i/_0829_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_2052_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/_0862_ ),
    .C1(\i_ibex/cs_registers_i/_0863_ ),
    .B1(\i_ibex/cs_registers_i/_0861_ ),
    .A1(net619),
    .Y(\i_ibex/cs_registers_i/_0864_ ),
    .A2(\i_ibex/cs_registers_i/_0833_ ));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2054_  (.Y(\i_ibex/cs_registers_i/_0866_ ),
    .A(net445),
    .B(net926),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout958 (.A(\i_ibex/cs_registers_i/csr_wdata_int [13]),
    .X(net958),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2056_  (.A(\i_ibex/cs_registers_i/dcsr_q [31]),
    .B(net909),
    .X(\i_ibex/cs_registers_i/dcsr_d [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2057_  (.Y(\i_ibex/cs_registers_i/dcsr_d [30]),
    .B(net908),
    .A_N(\i_ibex/cs_registers_i/dcsr_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2058_  (.A(\i_ibex/cs_registers_i/dcsr_q [21]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2059_  (.A(\i_ibex/cs_registers_i/dcsr_q [20]),
    .B(net909),
    .X(\i_ibex/cs_registers_i/dcsr_d [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2060_  (.A(\i_ibex/cs_registers_i/dcsr_q [19]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2061_  (.A(\i_ibex/cs_registers_i/dcsr_q [18]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2062_  (.A(\i_ibex/cs_registers_i/dcsr_q [17]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2063_  (.A(\i_ibex/cs_registers_i/dcsr_q [16]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/cs_registers_i/_2064_  (.A(net445),
    .B(net926),
    .X(\i_ibex/cs_registers_i/_0868_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2066_  (.A0(\i_ibex/debug_ebreakm ),
    .A1(net960),
    .S(\i_ibex/cs_registers_i/_0868_ ),
    .X(\i_ibex/cs_registers_i/dcsr_d [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2067_  (.A(\i_ibex/cs_registers_i/dcsr_q [14]),
    .B(net907),
    .X(\i_ibex/cs_registers_i/dcsr_d [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2068_  (.A0(\i_ibex/cs_registers_i/dcsr_q [13]),
    .A1(net957),
    .S(\i_ibex/cs_registers_i/_0868_ ),
    .X(\i_ibex/cs_registers_i/dcsr_d [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2069_  (.A(\i_ibex/debug_ebreaku ),
    .B(\i_ibex/cs_registers_i/_0868_ ),
    .Y(\i_ibex/cs_registers_i/_0870_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2070_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0548_ ),
    .A2(\i_ibex/cs_registers_i/_0868_ ),
    .Y(\i_ibex/cs_registers_i/dcsr_d [12]),
    .B1(\i_ibex/cs_registers_i/_0870_ ));
 sg13g2_buf_2 fanout956 (.A(\i_ibex/cs_registers_i/csr_wdata_int [7]),
    .X(net956),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2072_  (.A(\i_ibex/cs_registers_i/dcsr_q [29]),
    .B(net910),
    .X(\i_ibex/cs_registers_i/dcsr_d [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2073_  (.A(\i_ibex/cs_registers_i/dcsr_q [11]),
    .B(net910),
    .X(\i_ibex/cs_registers_i/dcsr_d [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2074_  (.A(\i_ibex/cs_registers_i/dcsr_q [10]),
    .B(net907),
    .X(\i_ibex/cs_registers_i/dcsr_d [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2075_  (.A(\i_ibex/cs_registers_i/dcsr_q [9]),
    .B(net907),
    .X(\i_ibex/cs_registers_i/dcsr_d [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2076_  (.A(\i_ibex/cs_registers_i/dcsr_q [5]),
    .B(net910),
    .X(\i_ibex/cs_registers_i/dcsr_d [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2077_  (.A(\i_ibex/cs_registers_i/dcsr_q [4]),
    .B(net907),
    .X(\i_ibex/cs_registers_i/dcsr_d [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2078_  (.A(\i_ibex/cs_registers_i/dcsr_q [3]),
    .B(net907),
    .X(\i_ibex/cs_registers_i/dcsr_d [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2079_  (.A0(\i_ibex/debug_single_step ),
    .A1(net949),
    .S(\i_ibex/cs_registers_i/_0868_ ),
    .X(\i_ibex/cs_registers_i/dcsr_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout955 (.X(net955),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2081_  (.A(\i_ibex/debug_csr_save ),
    .B(\i_ibex/csr_save_cause ),
    .X(\i_ibex/cs_registers_i/_0873_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout954 (.A(\i_ibex/cs_registers_i/csr_wdata_int [4]),
    .X(net954),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2084_  (.A(\i_ibex/cs_registers_i/dcsr_q [1]),
    .B(\i_ibex/cs_registers_i/_0868_ ),
    .Y(\i_ibex/cs_registers_i/_0876_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2085_  (.A(net971),
    .B(net973),
    .C(net907),
    .Y(\i_ibex/cs_registers_i/_0877_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2086_  (.A(\i_ibex/cs_registers_i/_0876_ ),
    .B(\i_ibex/cs_registers_i/_0877_ ),
    .C(net495),
    .Y(\i_ibex/cs_registers_i/_0878_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2087_  (.A2(net495),
    .A1(net785),
    .B1(\i_ibex/cs_registers_i/_0878_ ),
    .X(\i_ibex/cs_registers_i/dcsr_d [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2088_  (.A(\i_ibex/cs_registers_i/dcsr_q [0]),
    .B(\i_ibex/cs_registers_i/_0868_ ),
    .Y(\i_ibex/cs_registers_i/_0879_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2089_  (.A(\i_ibex/cs_registers_i/_0877_ ),
    .B(net495),
    .C(\i_ibex/cs_registers_i/_0879_ ),
    .Y(\i_ibex/cs_registers_i/_0880_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2090_  (.A2(net495),
    .A1(net786),
    .B1(\i_ibex/cs_registers_i/_0880_ ),
    .X(\i_ibex/cs_registers_i/dcsr_d [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2091_  (.A0(\i_ibex/cs_registers_i/dcsr_q [8]),
    .A1(\i_ibex/debug_cause [2]),
    .S(net492),
    .X(\i_ibex/cs_registers_i/dcsr_d [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2092_  (.A(\i_ibex/cs_registers_i/dcsr_q [28]),
    .B(net909),
    .X(\i_ibex/cs_registers_i/dcsr_d [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2093_  (.A0(\i_ibex/cs_registers_i/dcsr_q [7]),
    .A1(\i_ibex/debug_cause [1]),
    .S(net492),
    .X(\i_ibex/cs_registers_i/dcsr_d [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2094_  (.A0(\i_ibex/cs_registers_i/dcsr_q [6]),
    .A1(\i_ibex/debug_cause [0]),
    .S(net491),
    .X(\i_ibex/cs_registers_i/dcsr_d [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2095_  (.A(\i_ibex/cs_registers_i/dcsr_q [27]),
    .B(net907),
    .X(\i_ibex/cs_registers_i/dcsr_d [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2096_  (.A(\i_ibex/cs_registers_i/dcsr_q [26]),
    .B(net909),
    .X(\i_ibex/cs_registers_i/dcsr_d [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2097_  (.A(\i_ibex/cs_registers_i/dcsr_q [25]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2098_  (.A(\i_ibex/cs_registers_i/dcsr_q [24]),
    .B(net908),
    .X(\i_ibex/cs_registers_i/dcsr_d [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2099_  (.A(\i_ibex/cs_registers_i/dcsr_q [23]),
    .B(net909),
    .X(\i_ibex/cs_registers_i/dcsr_d [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2100_  (.A(\i_ibex/cs_registers_i/dcsr_q [22]),
    .B(net909),
    .X(\i_ibex/cs_registers_i/dcsr_d [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2101_  (.Y(\i_ibex/cs_registers_i/_0881_ ),
    .A(\i_ibex/debug_csr_save ),
    .B(\i_ibex/csr_save_cause ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2102_  (.Y(\i_ibex/cs_registers_i/dcsr_en ),
    .A(net907),
    .B(net1113),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout952 (.X(net952),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(net952),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2105_  (.A0(\i_ibex/pc_id [31]),
    .A1(\i_ibex/pc_if [31]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0884_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2106_  (.A0(net422),
    .A1(\i_ibex/cs_registers_i/_0884_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2108_  (.A0(\i_ibex/pc_id [30]),
    .A1(\i_ibex/pc_if [30]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0886_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2109_  (.A0(net963),
    .A1(\i_ibex/cs_registers_i/_0886_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2110_  (.A0(\i_ibex/pc_id [21]),
    .A1(\i_ibex/pc_if [21]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0887_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2111_  (.A0(net962),
    .A1(\i_ibex/cs_registers_i/_0887_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2112_  (.A0(\i_ibex/pc_id [20]),
    .A1(\i_ibex/pc_if [20]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0888_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2113_  (.A0(net426),
    .A1(\i_ibex/cs_registers_i/_0888_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2114_  (.A0(\i_ibex/pc_id [19]),
    .A1(\i_ibex/pc_if [19]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0889_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(net950),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2116_  (.A0(net947),
    .A1(\i_ibex/cs_registers_i/_0889_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2117_  (.A0(\i_ibex/pc_id [18]),
    .A1(\i_ibex/pc_if [18]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0891_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2118_  (.A0(net945),
    .A1(\i_ibex/cs_registers_i/_0891_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2119_  (.A0(\i_ibex/pc_id [17]),
    .A1(\i_ibex/pc_if [17]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0892_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2120_  (.A0(net944),
    .A1(\i_ibex/cs_registers_i/_0892_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2122_  (.A0(\i_ibex/pc_id [16]),
    .A1(\i_ibex/pc_if [16]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0894_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2123_  (.A0(net941),
    .A1(\i_ibex/cs_registers_i/_0894_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2124_  (.A0(\i_ibex/pc_id [15]),
    .A1(\i_ibex/pc_if [15]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0895_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2125_  (.A0(net960),
    .A1(\i_ibex/cs_registers_i/_0895_ ),
    .S(net492),
    .X(\i_ibex/cs_registers_i/depc_d [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2126_  (.A0(\i_ibex/pc_id [14]),
    .A1(\i_ibex/pc_if [14]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0896_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2127_  (.A(net1113),
    .B(\i_ibex/cs_registers_i/_0896_ ),
    .Y(\i_ibex/cs_registers_i/_0897_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2128_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0506_ ),
    .A2(net1113),
    .Y(\i_ibex/cs_registers_i/depc_d [14]),
    .B1(\i_ibex/cs_registers_i/_0897_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2129_  (.A0(\i_ibex/pc_id [13]),
    .A1(\i_ibex/pc_if [13]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0898_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2130_  (.A0(net957),
    .A1(\i_ibex/cs_registers_i/_0898_ ),
    .S(net492),
    .X(\i_ibex/cs_registers_i/depc_d [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2131_  (.A0(\i_ibex/pc_id [12]),
    .A1(\i_ibex/pc_if [12]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0899_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2132_  (.A(net1113),
    .B(\i_ibex/cs_registers_i/_0899_ ),
    .Y(\i_ibex/cs_registers_i/_0900_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2133_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0548_ ),
    .A2(\i_ibex/cs_registers_i/_0881_ ),
    .Y(\i_ibex/cs_registers_i/depc_d [12]),
    .B1(\i_ibex/cs_registers_i/_0900_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2134_  (.A0(\i_ibex/pc_id [29]),
    .A1(\i_ibex/pc_if [29]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0901_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2135_  (.A0(net421),
    .A1(\i_ibex/cs_registers_i/_0901_ ),
    .S(net492),
    .X(\i_ibex/cs_registers_i/depc_d [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2136_  (.A0(\i_ibex/pc_id [11]),
    .A1(\i_ibex/pc_if [11]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0902_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2137_  (.A0(net937),
    .A1(\i_ibex/cs_registers_i/_0902_ ),
    .S(net492),
    .X(\i_ibex/cs_registers_i/depc_d [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2138_  (.A0(\i_ibex/pc_id [10]),
    .A1(\i_ibex/pc_if [10]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0903_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2139_  (.A0(net935),
    .A1(\i_ibex/cs_registers_i/_0903_ ),
    .S(net492),
    .X(\i_ibex/cs_registers_i/depc_d [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2140_  (.A0(\i_ibex/pc_id [9]),
    .A1(\i_ibex/pc_if [9]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0904_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2141_  (.A0(net933),
    .A1(\i_ibex/cs_registers_i/_0904_ ),
    .S(net492),
    .X(\i_ibex/cs_registers_i/depc_d [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2142_  (.A0(\i_ibex/pc_id [8]),
    .A1(\i_ibex/pc_if [8]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0905_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(net948),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2144_  (.A0(net931),
    .A1(\i_ibex/cs_registers_i/_0905_ ),
    .S(net494),
    .X(\i_ibex/cs_registers_i/depc_d [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2145_  (.A0(\i_ibex/pc_id [7]),
    .A1(\i_ibex/pc_if [7]),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0907_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2146_  (.A0(net955),
    .A1(\i_ibex/cs_registers_i/_0907_ ),
    .S(net494),
    .X(\i_ibex/cs_registers_i/depc_d [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2147_  (.A0(\i_ibex/pc_id [6]),
    .A1(\i_ibex/pc_if [6]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0908_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2148_  (.A(net1113),
    .B(\i_ibex/cs_registers_i/_0908_ ),
    .Y(\i_ibex/cs_registers_i/_0909_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2149_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0682_ ),
    .A2(net1113),
    .Y(\i_ibex/cs_registers_i/depc_d [6]),
    .B1(\i_ibex/cs_registers_i/_0909_ ));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2150_  (.A0(\i_ibex/pc_id [5]),
    .A1(\i_ibex/pc_if [5]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0910_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2151_  (.A(net1113),
    .B(\i_ibex/cs_registers_i/_0910_ ),
    .Y(\i_ibex/cs_registers_i/_0911_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2152_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0195_ ),
    .A2(net1113),
    .Y(\i_ibex/cs_registers_i/depc_d [5]),
    .B1(\i_ibex/cs_registers_i/_0911_ ));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2153_  (.A0(\i_ibex/pc_id [4]),
    .A1(\i_ibex/pc_if [4]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0912_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2154_  (.A0(net953),
    .A1(\i_ibex/cs_registers_i/_0912_ ),
    .S(net494),
    .X(\i_ibex/cs_registers_i/depc_d [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2155_  (.A0(\i_ibex/pc_id [3]),
    .A1(\i_ibex/pc_if [3]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0913_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2156_  (.A0(net951),
    .A1(\i_ibex/cs_registers_i/_0913_ ),
    .S(net494),
    .X(\i_ibex/cs_registers_i/depc_d [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2157_  (.A0(\i_ibex/pc_id [2]),
    .A1(\i_ibex/pc_if [2]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0914_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2158_  (.A0(net950),
    .A1(\i_ibex/cs_registers_i/_0914_ ),
    .S(net494),
    .X(\i_ibex/cs_registers_i/depc_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2159_  (.A0(\i_ibex/pc_id [28]),
    .A1(\i_ibex/pc_if [28]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0915_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2160_  (.A0(net418),
    .A1(\i_ibex/cs_registers_i/_0915_ ),
    .S(net494),
    .X(\i_ibex/cs_registers_i/depc_d [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2161_  (.A0(\i_ibex/pc_id [1]),
    .A1(net1478),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0916_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2162_  (.A0(net971),
    .A1(\i_ibex/cs_registers_i/_0916_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2163_  (.A0(\i_ibex/pc_id [0]),
    .A1(net378),
    .S(net607),
    .X(\i_ibex/cs_registers_i/_0917_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2164_  (.A(net494),
    .B(\i_ibex/cs_registers_i/_0917_ ),
    .X(\i_ibex/cs_registers_i/depc_d [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2165_  (.A0(\i_ibex/pc_id [27]),
    .A1(\i_ibex/pc_if [27]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0918_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2166_  (.A0(net425),
    .A1(\i_ibex/cs_registers_i/_0918_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/cs_registers_i/_2167_  (.A0(\i_ibex/pc_id [26]),
    .A1(\i_ibex/pc_if [26]),
    .S(net609),
    .X(\i_ibex/cs_registers_i/_0919_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2168_  (.A0(net929),
    .A1(\i_ibex/cs_registers_i/_0919_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2169_  (.A0(\i_ibex/pc_id [25]),
    .A1(\i_ibex/pc_if [25]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0920_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2170_  (.A0(net416),
    .A1(\i_ibex/cs_registers_i/_0920_ ),
    .S(net493),
    .X(\i_ibex/cs_registers_i/depc_d [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2171_  (.A0(\i_ibex/pc_id [24]),
    .A1(\i_ibex/pc_if [24]),
    .S(net608),
    .X(\i_ibex/cs_registers_i/_0921_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2172_  (.A0(net927),
    .A1(\i_ibex/cs_registers_i/_0921_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2173_  (.A0(\i_ibex/pc_id [23]),
    .A1(\i_ibex/pc_if [23]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0922_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2174_  (.A0(net414),
    .A1(\i_ibex/cs_registers_i/_0922_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2175_  (.A0(\i_ibex/pc_id [22]),
    .A1(\i_ibex/pc_if [22]),
    .S(net606),
    .X(\i_ibex/cs_registers_i/_0923_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2176_  (.A0(net412),
    .A1(\i_ibex/cs_registers_i/_0923_ ),
    .S(net491),
    .X(\i_ibex/cs_registers_i/depc_d [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2177_  (.Y(\i_ibex/cs_registers_i/_0924_ ),
    .B1(\i_ibex/cs_registers_i/_0861_ ),
    .B2(\i_ibex/cs_registers_i/_0862_ ),
    .A2(\i_ibex/cs_registers_i/_0833_ ),
    .A1(net619),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/cs_registers_i/_2178_  (.Y(\i_ibex/cs_registers_i/_0925_ ),
    .B(\i_ibex/cs_registers_i/_0924_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/cs_registers_i/_0863_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2179_  (.Y(\i_ibex/cs_registers_i/_0926_ ),
    .A(\i_ibex/cs_registers_i/_0127_ ),
    .B(\i_ibex/cs_registers_i/_0286_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2180_  (.B1(\i_ibex/cs_registers_i/_0881_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/depc_en ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0925_ ),
    .A2(\i_ibex/cs_registers_i/_0926_ ));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2181_  (.Y(\i_ibex/cs_registers_i/_0927_ ),
    .A(\i_ibex/cs_registers_i/_0135_ ),
    .B(\i_ibex/cs_registers_i/_0864_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_2182_  (.A(net1094),
    .B(\i_ibex/cs_registers_i/_0056_ ),
    .C(\i_ibex/cs_registers_i/_0062_ ),
    .Y(\i_ibex/cs_registers_i/dscratch0_en ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_0927_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2183_  (.A(net450),
    .B(net926),
    .X(\i_ibex/cs_registers_i/dscratch1_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2184_  (.Y(\i_ibex/cs_registers_i/_0928_ ),
    .A(net784),
    .B(net926),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_2185_  (.A(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_q ),
    .B(\i_ibex/cs_registers_i/_0081_ ),
    .C(\i_ibex/cs_registers_i/_0329_ ),
    .D(\i_ibex/cs_registers_i/_0928_ ),
    .Y(\i_ibex/cs_registers_i/gen_trigger_regs.tmatch_control_we ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2186_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0929_ ),
    .A(net446),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2187_  (.A(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_q ),
    .B(\i_ibex/cs_registers_i/_0929_ ),
    .C(\i_ibex/cs_registers_i/_0928_ ),
    .Y(\i_ibex/cs_registers_i/gen_trigger_regs.tmatch_value_we ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2188_  (.A(\i_ibex/cs_registers_i/_0027_ ),
    .B(\i_ibex/cs_registers_i/_0329_ ),
    .C(\i_ibex/cs_registers_i/_0928_ ),
    .Y(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_we ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 \i_ibex/cs_registers_i/_2189_  (.A(\i_ibex/cs_registers_i/_0924_ ),
    .Y(\i_ibex/illegal_csr_insn_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2190_  (.A(\i_ibex/perf_instr_ret_wb ),
    .B(\i_ibex/cs_registers_i/instr_ret_i_$_AND__A_B ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i_counter_inc_i ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2191_  (.A(irqs_i[7]),
    .B(\i_ibex/cs_registers_i/mie_q [7]),
    .X(\i_ibex/irqs [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2192_  (.A(net35),
    .B(\i_ibex/cs_registers_i/mie_q [18]),
    .X(\i_ibex/irqs [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2193_  (.A(irqs_i[9]),
    .B(\i_ibex/cs_registers_i/mie_q [9]),
    .X(\i_ibex/irqs [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2194_  (.A(\i_ibex/irqs [7]),
    .B(\i_ibex/irqs [18]),
    .C(\i_ibex/irqs [9]),
    .Y(\i_ibex/cs_registers_i/_0930_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2195_  (.A(irqs_i[3]),
    .B(\i_ibex/cs_registers_i/mie_q [3]),
    .X(\i_ibex/irqs [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2196_  (.A(timer0_irq_i),
    .B(\i_ibex/cs_registers_i/mie_q [17]),
    .X(\i_ibex/irqs [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2197_  (.A(\i_ibex/irqs [3]),
    .B(\i_ibex/irqs [17]),
    .Y(\i_ibex/cs_registers_i/_0931_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2198_  (.A(irqs_i[4]),
    .B(\i_ibex/cs_registers_i/mie_q [4]),
    .X(\i_ibex/irqs [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2199_  (.A(irqs_i[5]),
    .B(\i_ibex/cs_registers_i/mie_q [5]),
    .X(\i_ibex/irqs [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2200_  (.A(\i_ibex/irqs [4]),
    .B(\i_ibex/irqs [5]),
    .Y(\i_ibex/cs_registers_i/_0932_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2201_  (.A(irqs_i[6]),
    .B(\i_ibex/cs_registers_i/mie_q [6]),
    .X(\i_ibex/irqs [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2202_  (.A(irqs_i[0]),
    .B(\i_ibex/cs_registers_i/mie_q [0]),
    .X(\i_ibex/irqs [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2203_  (.A(\i_ibex/irqs [6]),
    .B(\i_ibex/irqs [0]),
    .Y(\i_ibex/cs_registers_i/_0933_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2204_  (.A(irqs_i[8]),
    .B(\i_ibex/cs_registers_i/mie_q [8]),
    .X(\i_ibex/irqs [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2205_  (.A(irqs_i[1]),
    .B(\i_ibex/cs_registers_i/mie_q [1]),
    .X(\i_ibex/irqs [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2206_  (.A(\i_ibex/irqs [8]),
    .B(\i_ibex/irqs [1]),
    .Y(\i_ibex/cs_registers_i/_0934_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/_2207_  (.A(\i_ibex/cs_registers_i/_0931_ ),
    .B(\i_ibex/cs_registers_i/_0932_ ),
    .C(\i_ibex/cs_registers_i/_0933_ ),
    .D(\i_ibex/cs_registers_i/_0934_ ),
    .X(\i_ibex/cs_registers_i/_0935_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2208_  (.A(irqs_i[2]),
    .B(\i_ibex/cs_registers_i/mie_q [2]),
    .X(\i_ibex/irqs [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2209_  (.A(irqs_i[10]),
    .B(\i_ibex/cs_registers_i/mie_q [10]),
    .X(\i_ibex/irqs [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2210_  (.A(\i_ibex/irqs [2]),
    .B(\i_ibex/irqs [10]),
    .Y(\i_ibex/cs_registers_i/_0936_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2211_  (.A(irqs_i[15]),
    .B(\i_ibex/cs_registers_i/mie_q [15]),
    .X(\i_ibex/irqs [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2212_  (.A(net36),
    .B(\i_ibex/cs_registers_i/mie_q [16]),
    .X(\i_ibex/irqs [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2213_  (.A(\i_ibex/irqs [15]),
    .B(\i_ibex/irqs [16]),
    .Y(\i_ibex/cs_registers_i/_0937_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2214_  (.A(irqs_i[11]),
    .B(\i_ibex/cs_registers_i/mie_q [11]),
    .X(\i_ibex/irqs [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2215_  (.A(irqs_i[12]),
    .B(\i_ibex/cs_registers_i/mie_q [12]),
    .X(\i_ibex/irqs [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2216_  (.A(\i_ibex/irqs [11]),
    .B(\i_ibex/irqs [12]),
    .Y(\i_ibex/cs_registers_i/_0938_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2217_  (.A(irqs_i[13]),
    .B(\i_ibex/cs_registers_i/mie_q [13]),
    .X(\i_ibex/irqs [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2218_  (.A(irqs_i[14]),
    .B(\i_ibex/cs_registers_i/mie_q [14]),
    .X(\i_ibex/irqs [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2219_  (.A(\i_ibex/irqs [13]),
    .B(\i_ibex/irqs [14]),
    .Y(\i_ibex/cs_registers_i/_0939_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/_2220_  (.A(\i_ibex/cs_registers_i/_0936_ ),
    .B(\i_ibex/cs_registers_i/_0937_ ),
    .C(\i_ibex/cs_registers_i/_0938_ ),
    .D(\i_ibex/cs_registers_i/_0939_ ),
    .X(\i_ibex/cs_registers_i/_0940_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2221_  (.B(\i_ibex/cs_registers_i/_0935_ ),
    .C(\i_ibex/cs_registers_i/_0940_ ),
    .A(\i_ibex/cs_registers_i/_0930_ ),
    .Y(\i_ibex/irq_pending_o ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_2222_  (.A(\i_ibex/debug_csr_save ),
    .B_N(\i_ibex/csr_save_cause ),
    .Y(\i_ibex/cs_registers_i/_0941_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2223_  (.Y(\i_ibex/cs_registers_i/_0942_ ),
    .A(\i_ibex/cs_registers_i/_0831_ ),
    .B(\i_ibex/cs_registers_i/_0941_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/cs_registers_i/_2224_  (.Y(\i_ibex/cs_registers_i/_0943_ ),
    .B(net624),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/csr_save_cause ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2225_  (.A(net480),
    .B(\i_ibex/cs_registers_i/_0943_ ),
    .X(\i_ibex/cs_registers_i/_0944_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2226_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0945_ ),
    .A(\i_ibex/cs_registers_i/_0944_ ),
    .VSS(VSS));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2228_  (.Y(\i_ibex/cs_registers_i/_0947_ ),
    .B(\i_ibex/csr_restore_mret_id ),
    .A_N(\i_ibex/nmi_mode ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2229_  (.Y(\i_ibex/cs_registers_i/_0948_ ),
    .A(\i_ibex/cs_registers_i/_0945_ ),
    .B(\i_ibex/cs_registers_i/_0947_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout945 (.X(net945),
    .A(net946),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/cs_registers_i/_2231_  (.A(net624),
    .B(\i_ibex/nmi_mode ),
    .X(\i_ibex/cs_registers_i/_0950_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_16 \i_ibex/cs_registers_i/_2233_  (.A(\i_ibex/cs_registers_i/_0942_ ),
    .Y(\i_ibex/cs_registers_i/_0952_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2235_  (.Y(\i_ibex/cs_registers_i/_0954_ ),
    .B1(net1057),
    .B2(\i_ibex/exc_cause [6]),
    .A2(net1268),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2236_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0955_ ),
    .A(\i_ibex/cs_registers_i/_0954_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2237_  (.A2(net1022),
    .A1(net423),
    .B1(\i_ibex/cs_registers_i/_0955_ ),
    .X(\i_ibex/cs_registers_i/mcause_d [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/_2238_  (.A(\i_ibex/cs_registers_i/_0944_ ),
    .B_N(\i_ibex/cs_registers_i/_0947_ ),
    .Y(\i_ibex/cs_registers_i/_0956_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(net942),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2241_  (.Y(\i_ibex/cs_registers_i/_0959_ ),
    .B1(net1055),
    .B2(\i_ibex/exc_cause [5]),
    .A2(net1267),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2242_  (.B1(\i_ibex/cs_registers_i/_0959_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcause_d [5]),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0195_ ),
    .A2(\i_ibex/cs_registers_i/_0956_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2243_  (.Y(\i_ibex/cs_registers_i/_0960_ ),
    .B1(net1053),
    .B2(\i_ibex/exc_cause [4]),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2244_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0961_ ),
    .A(\i_ibex/cs_registers_i/_0960_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2245_  (.A2(net1022),
    .A1(net953),
    .B1(\i_ibex/cs_registers_i/_0961_ ),
    .X(\i_ibex/cs_registers_i/mcause_d [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_2246_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_0962_ ),
    .B(\i_ibex/csr_save_cause ),
    .A(\i_ibex/csr_restore_mret_id ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2247_  (.B1(\i_ibex/csr_save_cause ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0963_ ),
    .VSS(VSS),
    .A1(net784),
    .A2(\i_ibex/debug_csr_save ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2248_  (.B(\i_ibex/cs_registers_i/_0962_ ),
    .C(\i_ibex/cs_registers_i/_0963_ ),
    .A(\i_ibex/cs_registers_i/_0947_ ),
    .Y(\i_ibex/cs_registers_i/_0964_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2249_  (.Y(\i_ibex/cs_registers_i/_0965_ ),
    .A(net951),
    .B(\i_ibex/cs_registers_i/_0964_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2252_  (.Y(\i_ibex/cs_registers_i/_0967_ ),
    .B1(net1053),
    .B2(\i_ibex/exc_cause [3]),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2253_  (.Y(\i_ibex/cs_registers_i/mcause_d [3]),
    .A(\i_ibex/cs_registers_i/_0965_ ),
    .B(\i_ibex/cs_registers_i/_0967_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2254_  (.Y(\i_ibex/cs_registers_i/_0968_ ),
    .B1(net1053),
    .B2(\i_ibex/exc_cause [2]),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2255_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0969_ ),
    .A(\i_ibex/cs_registers_i/_0968_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2256_  (.A2(\i_ibex/cs_registers_i/_0964_ ),
    .A1(net950),
    .B1(\i_ibex/cs_registers_i/_0969_ ),
    .X(\i_ibex/cs_registers_i/mcause_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2257_  (.Y(\i_ibex/cs_registers_i/_0970_ ),
    .A(net971),
    .B(\i_ibex/cs_registers_i/_0964_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2258_  (.Y(\i_ibex/cs_registers_i/_0971_ ),
    .B1(net1054),
    .B2(\i_ibex/exc_cause [1]),
    .A2(net1266),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2259_  (.Y(\i_ibex/cs_registers_i/mcause_d [1]),
    .A(\i_ibex/cs_registers_i/_0970_ ),
    .B(\i_ibex/cs_registers_i/_0971_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2260_  (.Y(\i_ibex/cs_registers_i/_0972_ ),
    .A(net973),
    .B(\i_ibex/cs_registers_i/_0964_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2261_  (.Y(\i_ibex/cs_registers_i/_0973_ ),
    .B1(net1054),
    .B2(\i_ibex/exc_cause [0]),
    .A2(net1266),
    .A1(\i_ibex/cs_registers_i/mstack_cause_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2262_  (.Y(\i_ibex/cs_registers_i/mcause_d [0]),
    .A(\i_ibex/cs_registers_i/_0972_ ),
    .B(\i_ibex/cs_registers_i/_0973_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2263_  (.A(net1268),
    .B(net1057),
    .Y(\i_ibex/cs_registers_i/_0974_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2264_  (.B1(\i_ibex/cs_registers_i/_0974_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcause_en ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0072_ ),
    .A2(\i_ibex/cs_registers_i/_0927_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2265_  (.Y(\i_ibex/cs_registers_i/_0975_ ),
    .A(net983),
    .B(net926),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2266_  (.A0(net973),
    .A1(\i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y [192]),
    .S(\i_ibex/cs_registers_i/_0975_ ),
    .X(\i_ibex/cs_registers_i/_0002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2267_  (.A0(net949),
    .A1(\i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y [194]),
    .S(\i_ibex/cs_registers_i/_0975_ ),
    .X(\i_ibex/cs_registers_i/_0003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2268_  (.Y(\i_ibex/cs_registers_i/_0976_ ),
    .B1(net1059),
    .B2(\i_ibex/cs_registers_i/_0884_ ),
    .A2(net1270),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2269_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0977_ ),
    .A(\i_ibex/cs_registers_i/_0976_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2270_  (.A2(net1020),
    .A1(net423),
    .B1(\i_ibex/cs_registers_i/_0977_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout938 (.A(\i_ibex/cs_registers_i/csr_wdata_int [11]),
    .X(net938),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2272_  (.Y(\i_ibex/cs_registers_i/_0979_ ),
    .A(net963),
    .B(net1020),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2273_  (.Y(\i_ibex/cs_registers_i/_0980_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0886_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2274_  (.Y(\i_ibex/cs_registers_i/mepc_d [30]),
    .A(\i_ibex/cs_registers_i/_0979_ ),
    .B(\i_ibex/cs_registers_i/_0980_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2275_  (.Y(\i_ibex/cs_registers_i/_0981_ ),
    .A(net962),
    .B(net1020),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2276_  (.Y(\i_ibex/cs_registers_i/_0982_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0887_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2277_  (.Y(\i_ibex/cs_registers_i/mepc_d [21]),
    .A(\i_ibex/cs_registers_i/_0981_ ),
    .B(\i_ibex/cs_registers_i/_0982_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2278_  (.Y(\i_ibex/cs_registers_i/_0983_ ),
    .A(net426),
    .B(net1019),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2279_  (.Y(\i_ibex/cs_registers_i/_0984_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0888_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2280_  (.Y(\i_ibex/cs_registers_i/mepc_d [20]),
    .A(\i_ibex/cs_registers_i/_0983_ ),
    .B(\i_ibex/cs_registers_i/_0984_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2282_  (.Y(\i_ibex/cs_registers_i/_0986_ ),
    .B1(net1059),
    .B2(\i_ibex/cs_registers_i/_0889_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2283_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0987_ ),
    .A(\i_ibex/cs_registers_i/_0986_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2284_  (.A2(net1019),
    .A1(net947),
    .B1(\i_ibex/cs_registers_i/_0987_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2285_  (.Y(\i_ibex/cs_registers_i/_0988_ ),
    .B1(net1059),
    .B2(\i_ibex/cs_registers_i/_0891_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2286_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0989_ ),
    .A(\i_ibex/cs_registers_i/_0988_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2287_  (.A2(net1019),
    .A1(net945),
    .B1(\i_ibex/cs_registers_i/_0989_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2288_  (.Y(\i_ibex/cs_registers_i/_0990_ ),
    .A(net944),
    .B(net1020),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2289_  (.Y(\i_ibex/cs_registers_i/_0991_ ),
    .B1(net1059),
    .B2(\i_ibex/cs_registers_i/_0892_ ),
    .A2(net1270),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2290_  (.Y(\i_ibex/cs_registers_i/mepc_d [17]),
    .A(\i_ibex/cs_registers_i/_0990_ ),
    .B(\i_ibex/cs_registers_i/_0991_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout936 (.A(\i_ibex/cs_registers_i/csr_wdata_int [10]),
    .X(net936),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2292_  (.Y(\i_ibex/cs_registers_i/_0993_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0894_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2293_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_0994_ ),
    .A(\i_ibex/cs_registers_i/_0993_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2294_  (.A2(net1020),
    .A1(net941),
    .B1(\i_ibex/cs_registers_i/_0994_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2295_  (.Y(\i_ibex/cs_registers_i/_0995_ ),
    .A(net960),
    .B(net1021),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2296_  (.Y(\i_ibex/cs_registers_i/_0996_ ),
    .B1(net1060),
    .B2(\i_ibex/cs_registers_i/_0895_ ),
    .A2(net1271),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2297_  (.Y(\i_ibex/cs_registers_i/mepc_d [15]),
    .A(\i_ibex/cs_registers_i/_0995_ ),
    .B(\i_ibex/cs_registers_i/_0996_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2298_  (.Y(\i_ibex/cs_registers_i/_0997_ ),
    .B1(net1057),
    .B2(\i_ibex/cs_registers_i/_0896_ ),
    .A2(net1268),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2299_  (.B1(\i_ibex/cs_registers_i/_0997_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mepc_d [14]),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0506_ ),
    .A2(\i_ibex/cs_registers_i/_0956_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2300_  (.Y(\i_ibex/cs_registers_i/_0998_ ),
    .A(net957),
    .B(net1021),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2301_  (.Y(\i_ibex/cs_registers_i/_0999_ ),
    .B1(net1060),
    .B2(\i_ibex/cs_registers_i/_0898_ ),
    .A2(net1271),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2302_  (.Y(\i_ibex/cs_registers_i/mepc_d [13]),
    .A(\i_ibex/cs_registers_i/_0998_ ),
    .B(\i_ibex/cs_registers_i/_0999_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2303_  (.Y(\i_ibex/cs_registers_i/_1000_ ),
    .B1(net1057),
    .B2(\i_ibex/cs_registers_i/_0899_ ),
    .A2(net1268),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2304_  (.B1(\i_ibex/cs_registers_i/_1000_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mepc_d [12]),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0548_ ),
    .A2(\i_ibex/cs_registers_i/_0956_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2305_  (.Y(\i_ibex/cs_registers_i/_1001_ ),
    .A(net421),
    .B(net1021),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2306_  (.Y(\i_ibex/cs_registers_i/_1002_ ),
    .B1(net1060),
    .B2(\i_ibex/cs_registers_i/_0901_ ),
    .A2(net1271),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2307_  (.Y(\i_ibex/cs_registers_i/mepc_d [29]),
    .A(\i_ibex/cs_registers_i/_1001_ ),
    .B(\i_ibex/cs_registers_i/_1002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2308_  (.Y(\i_ibex/cs_registers_i/_1003_ ),
    .A(net938),
    .B(net1022),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2309_  (.Y(\i_ibex/cs_registers_i/_1004_ ),
    .B1(net1057),
    .B2(\i_ibex/cs_registers_i/_0902_ ),
    .A2(net1268),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2310_  (.Y(\i_ibex/cs_registers_i/mepc_d [11]),
    .A(\i_ibex/cs_registers_i/_1003_ ),
    .B(\i_ibex/cs_registers_i/_1004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2311_  (.Y(\i_ibex/cs_registers_i/_1005_ ),
    .B1(\i_ibex/cs_registers_i/_0952_ ),
    .B2(\i_ibex/cs_registers_i/_0903_ ),
    .A2(net1268),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2312_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1006_ ),
    .A(\i_ibex/cs_registers_i/_1005_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2313_  (.A2(net1022),
    .A1(net936),
    .B1(\i_ibex/cs_registers_i/_1006_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2314_  (.Y(\i_ibex/cs_registers_i/_1007_ ),
    .B1(net1057),
    .B2(\i_ibex/cs_registers_i/_0904_ ),
    .A2(net1268),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2315_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1008_ ),
    .A(\i_ibex/cs_registers_i/_1007_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2316_  (.A2(net1022),
    .A1(net934),
    .B1(\i_ibex/cs_registers_i/_1008_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2317_  (.Y(\i_ibex/cs_registers_i/_1009_ ),
    .B1(net1053),
    .B2(\i_ibex/cs_registers_i/_0905_ ),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2318_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1010_ ),
    .A(\i_ibex/cs_registers_i/_1009_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2319_  (.A2(net1022),
    .A1(net932),
    .B1(\i_ibex/cs_registers_i/_1010_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2320_  (.Y(\i_ibex/cs_registers_i/_1011_ ),
    .A(net955),
    .B(net1022),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2321_  (.Y(\i_ibex/cs_registers_i/_1012_ ),
    .B1(net1053),
    .B2(\i_ibex/cs_registers_i/_0907_ ),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2322_  (.Y(\i_ibex/cs_registers_i/mepc_d [7]),
    .A(\i_ibex/cs_registers_i/_1011_ ),
    .B(\i_ibex/cs_registers_i/_1012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2323_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1013_ ),
    .A(\i_ibex/cs_registers_i/_0964_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2324_  (.Y(\i_ibex/cs_registers_i/_1014_ ),
    .B1(net1055),
    .B2(\i_ibex/cs_registers_i/_0908_ ),
    .A2(net1267),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2325_  (.B1(\i_ibex/cs_registers_i/_1014_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mepc_d [6]),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0682_ ),
    .A2(\i_ibex/cs_registers_i/_1013_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2326_  (.Y(\i_ibex/cs_registers_i/_1015_ ),
    .B1(net1055),
    .B2(\i_ibex/cs_registers_i/_0910_ ),
    .A2(net1267),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2327_  (.B1(\i_ibex/cs_registers_i/_1015_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mepc_d [5]),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0195_ ),
    .A2(\i_ibex/cs_registers_i/_1013_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2328_  (.Y(\i_ibex/cs_registers_i/_1016_ ),
    .B1(net1054),
    .B2(\i_ibex/cs_registers_i/_0912_ ),
    .A2(net1266),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2329_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1017_ ),
    .A(\i_ibex/cs_registers_i/_1016_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2330_  (.A2(net1022),
    .A1(net953),
    .B1(\i_ibex/cs_registers_i/_1017_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2331_  (.Y(\i_ibex/cs_registers_i/_1018_ ),
    .B1(net1053),
    .B2(\i_ibex/cs_registers_i/_0913_ ),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2332_  (.Y(\i_ibex/cs_registers_i/mepc_d [3]),
    .A(\i_ibex/cs_registers_i/_0965_ ),
    .B(\i_ibex/cs_registers_i/_1018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2333_  (.Y(\i_ibex/cs_registers_i/_1019_ ),
    .B1(net1054),
    .B2(\i_ibex/cs_registers_i/_0914_ ),
    .A2(net1266),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2334_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1020_ ),
    .A(\i_ibex/cs_registers_i/_1019_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2335_  (.A2(\i_ibex/cs_registers_i/_0964_ ),
    .A1(net950),
    .B1(\i_ibex/cs_registers_i/_1020_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2336_  (.Y(\i_ibex/cs_registers_i/_1021_ ),
    .B1(net1060),
    .B2(\i_ibex/cs_registers_i/_0915_ ),
    .A2(net1271),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2337_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1022_ ),
    .A(\i_ibex/cs_registers_i/_1021_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2338_  (.A2(net1021),
    .A1(net419),
    .B1(\i_ibex/cs_registers_i/_1022_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2339_  (.Y(\i_ibex/cs_registers_i/_1023_ ),
    .B1(net1053),
    .B2(\i_ibex/cs_registers_i/_0916_ ),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2340_  (.Y(\i_ibex/cs_registers_i/mepc_d [1]),
    .A(\i_ibex/cs_registers_i/_0970_ ),
    .B(\i_ibex/cs_registers_i/_1023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2341_  (.Y(\i_ibex/cs_registers_i/_1024_ ),
    .B1(net1053),
    .B2(\i_ibex/cs_registers_i/_0917_ ),
    .A2(net1265),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2342_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mepc_d [0]),
    .A(\i_ibex/cs_registers_i/_1024_ ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2343_  (.Y(\i_ibex/cs_registers_i/_1025_ ),
    .A(net425),
    .B(net1021),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2344_  (.Y(\i_ibex/cs_registers_i/_1026_ ),
    .B1(net1060),
    .B2(\i_ibex/cs_registers_i/_0918_ ),
    .A2(net1271),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2345_  (.Y(\i_ibex/cs_registers_i/mepc_d [27]),
    .A(\i_ibex/cs_registers_i/_1025_ ),
    .B(\i_ibex/cs_registers_i/_1026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2346_  (.Y(\i_ibex/cs_registers_i/_1027_ ),
    .B1(net1059),
    .B2(\i_ibex/cs_registers_i/_0919_ ),
    .A2(net1270),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2347_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1028_ ),
    .A(\i_ibex/cs_registers_i/_1027_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2348_  (.A2(net1019),
    .A1(net929),
    .B1(\i_ibex/cs_registers_i/_1028_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2349_  (.Y(\i_ibex/cs_registers_i/_1029_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0920_ ),
    .A2(net1270),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2350_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1030_ ),
    .A(\i_ibex/cs_registers_i/_1029_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2351_  (.A2(net1019),
    .A1(net417),
    .B1(\i_ibex/cs_registers_i/_1030_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2352_  (.Y(\i_ibex/cs_registers_i/_1031_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0921_ ),
    .A2(net1270),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2353_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1032_ ),
    .A(\i_ibex/cs_registers_i/_1031_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2354_  (.A2(net1019),
    .A1(net927),
    .B1(\i_ibex/cs_registers_i/_1032_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2355_  (.Y(\i_ibex/cs_registers_i/_1033_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0922_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2356_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1034_ ),
    .A(\i_ibex/cs_registers_i/_1033_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2357_  (.A2(net1019),
    .A1(net415),
    .B1(\i_ibex/cs_registers_i/_1034_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2358_  (.Y(\i_ibex/cs_registers_i/_1035_ ),
    .B1(net1058),
    .B2(\i_ibex/cs_registers_i/_0923_ ),
    .A2(net1269),
    .A1(\i_ibex/cs_registers_i/mstack_epc_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2359_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1036_ ),
    .A(\i_ibex/cs_registers_i/_1035_ ),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2360_  (.A2(net1019),
    .A1(net413),
    .B1(\i_ibex/cs_registers_i/_1036_ ),
    .X(\i_ibex/cs_registers_i/mepc_d [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2361_  (.Y(\i_ibex/cs_registers_i/_1037_ ),
    .A(net455),
    .B(net926),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2362_  (.B1(\i_ibex/cs_registers_i/_0974_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mepc_en ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0081_ ),
    .A2(\i_ibex/cs_registers_i/_1037_ ));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2363_  (.Y(\i_ibex/cs_registers_i/_1038_ ),
    .A(\i_ibex/cs_registers_i/_0081_ ),
    .B(\i_ibex/cs_registers_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_2364_  (.A(\i_ibex/cs_registers_i/_0103_ ),
    .B(\i_ibex/cs_registers_i/_0927_ ),
    .C(\i_ibex/cs_registers_i/_1038_ ),
    .Y(\i_ibex/cs_registers_i/mhpmcounter_we [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_2365_  (.A(\i_ibex/cs_registers_i/_0118_ ),
    .B(\i_ibex/cs_registers_i/_0925_ ),
    .C(\i_ibex/cs_registers_i/_1038_ ),
    .Y(\i_ibex/cs_registers_i/mhpmcounter_we [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/_2366_  (.A(\i_ibex/cs_registers_i/_0107_ ),
    .B(\i_ibex/cs_registers_i/_0927_ ),
    .C(\i_ibex/cs_registers_i/_1038_ ),
    .Y(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_2367_  (.A(\i_ibex/cs_registers_i/_0027_ ),
    .B(\i_ibex/cs_registers_i/_0107_ ),
    .C(\i_ibex/cs_registers_i/_0925_ ),
    .Y(\i_ibex/cs_registers_i/mhpmcounterh_we [0]),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1038_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2368_  (.A(net436),
    .B(net926),
    .X(\i_ibex/cs_registers_i/mie_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2369_  (.A(\i_ibex/cs_registers_i/_0027_ ),
    .B(\i_ibex/cs_registers_i/_1037_ ),
    .Y(\i_ibex/cs_registers_i/mscratch_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2370_  (.A(\i_ibex/cs_registers_i/_0027_ ),
    .B(\i_ibex/cs_registers_i/_0370_ ),
    .C(\i_ibex/cs_registers_i/_0863_ ),
    .Y(\i_ibex/cs_registers_i/_1039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/_2371_  (.Y(\i_ibex/cs_registers_i/_1040_ ),
    .A(\i_ibex/cs_registers_i/_0924_ ),
    .B(\i_ibex/cs_registers_i/_1039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2372_  (.A0(net951),
    .A1(\i_ibex/csr_mstatus_mie ),
    .S(net911),
    .X(\i_ibex/cs_registers_i/_1041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/_2373_  (.A(net624),
    .B(\i_ibex/cs_registers_i/mstatus_q [4]),
    .X(\i_ibex/cs_registers_i/_1042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/_2374_  (.A2(\i_ibex/cs_registers_i/_1041_ ),
    .A1(\i_ibex/cs_registers_i/_0944_ ),
    .B1(\i_ibex/cs_registers_i/_1042_ ),
    .X(\i_ibex/cs_registers_i/mstatus_d [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2375_  (.Y(\i_ibex/cs_registers_i/_1043_ ),
    .B(net911),
    .A_N(\i_ibex/cs_registers_i/mstatus_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2376_  (.B1(\i_ibex/cs_registers_i/_1043_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1044_ ),
    .VSS(VSS),
    .A1(net956),
    .A2(net911));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2377_  (.Y(\i_ibex/cs_registers_i/_1045_ ),
    .B(\i_ibex/nmi_mode ),
    .A_N(\i_ibex/cs_registers_i/mstack_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2378_  (.Y(\i_ibex/cs_registers_i/_1046_ ),
    .B1(\i_ibex/cs_registers_i/_1045_ ),
    .B2(\i_ibex/csr_restore_mret_id ),
    .A2(net1055),
    .A1(\i_ibex/csr_mstatus_mie ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2379_  (.B1(\i_ibex/cs_registers_i/_1046_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mstatus_d [4]),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0945_ ),
    .A2(\i_ibex/cs_registers_i/_1044_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/_2380_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/_1047_ ),
    .B(net559),
    .A(net564));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2381_  (.B1(\i_ibex/cs_registers_i/_0593_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1048_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_rdata [11]),
    .A2(\i_ibex/cs_registers_i/_1047_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2382_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1049_ ),
    .A(net559),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2383_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_1049_ ),
    .A2(\i_ibex/csr_rdata [11]),
    .Y(\i_ibex/cs_registers_i/_1050_ ),
    .B1(net631));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2384_  (.A(net564),
    .B(net559),
    .C(net691),
    .Y(\i_ibex/cs_registers_i/_1051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_2385_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net564),
    .C1(\i_ibex/cs_registers_i/_1051_ ),
    .B1(\i_ibex/cs_registers_i/_1050_ ),
    .A1(\i_ibex/cs_registers_i/_0546_ ),
    .Y(\i_ibex/cs_registers_i/_1052_ ),
    .A2(\i_ibex/cs_registers_i/_1048_ ));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2386_  (.Y(\i_ibex/cs_registers_i/_1053_ ),
    .B(net1055),
    .A_N(net785),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2387_  (.Y(\i_ibex/cs_registers_i/_1054_ ),
    .A(\i_ibex/cs_registers_i/_0943_ ),
    .B(\i_ibex/cs_registers_i/_1053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2388_  (.A0(net785),
    .A1(\i_ibex/cs_registers_i/mstatus_q [3]),
    .S(net784),
    .X(\i_ibex/cs_registers_i/_1055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2389_  (.Y(\i_ibex/cs_registers_i/_1056_ ),
    .A(\i_ibex/cs_registers_i/_0941_ ),
    .B(\i_ibex/cs_registers_i/_1055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2390_  (.B1(\i_ibex/cs_registers_i/_1056_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1057_ ),
    .VSS(VSS),
    .A1(net911),
    .A2(\i_ibex/cs_registers_i/_1054_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2391_  (.Y(\i_ibex/cs_registers_i/_1058_ ),
    .A(\i_ibex/cs_registers_i/_1052_ ),
    .B(\i_ibex/cs_registers_i/_1057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2392_  (.B(\i_ibex/cs_registers_i/_0943_ ),
    .C(net911),
    .A(\i_ibex/cs_registers_i/mstatus_q [3]),
    .Y(\i_ibex/cs_registers_i/_1059_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1053_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2393_  (.Y(\i_ibex/cs_registers_i/_1060_ ),
    .B1(net1055),
    .B2(net785),
    .A2(net1267),
    .A1(\i_ibex/cs_registers_i/mstack_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2394_  (.B(\i_ibex/cs_registers_i/_1059_ ),
    .C(\i_ibex/cs_registers_i/_1060_ ),
    .A(\i_ibex/cs_registers_i/_1058_ ),
    .Y(\i_ibex/cs_registers_i/mstatus_d [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/_2395_  (.Y(\i_ibex/cs_registers_i/_1061_ ),
    .B(net1055),
    .A_N(net786),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2396_  (.Y(\i_ibex/cs_registers_i/_1062_ ),
    .A(\i_ibex/cs_registers_i/_0943_ ),
    .B(\i_ibex/cs_registers_i/_1061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2397_  (.A0(net786),
    .A1(\i_ibex/cs_registers_i/mstatus_q [2]),
    .S(net784),
    .X(\i_ibex/cs_registers_i/_1063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2398_  (.Y(\i_ibex/cs_registers_i/_1064_ ),
    .A(\i_ibex/cs_registers_i/_0941_ ),
    .B(\i_ibex/cs_registers_i/_1063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2399_  (.B1(\i_ibex/cs_registers_i/_1064_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1065_ ),
    .VSS(VSS),
    .A1(net911),
    .A2(\i_ibex/cs_registers_i/_1062_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/_2400_  (.Y(\i_ibex/cs_registers_i/_1066_ ),
    .A(\i_ibex/cs_registers_i/_1052_ ),
    .B(\i_ibex/cs_registers_i/_1065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2401_  (.B(\i_ibex/cs_registers_i/_0943_ ),
    .C(net911),
    .A(\i_ibex/cs_registers_i/mstatus_q [2]),
    .Y(\i_ibex/cs_registers_i/_1067_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1061_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/_2402_  (.Y(\i_ibex/cs_registers_i/_1068_ ),
    .B1(net1055),
    .B2(net786),
    .A2(net1267),
    .A1(\i_ibex/cs_registers_i/mstack_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2403_  (.B(\i_ibex/cs_registers_i/_1067_ ),
    .C(\i_ibex/cs_registers_i/_1068_ ),
    .A(\i_ibex/cs_registers_i/_1066_ ),
    .Y(\i_ibex/cs_registers_i/mstatus_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2404_  (.A0(net961),
    .A1(\i_ibex/csr_mstatus_tw ),
    .S(\i_ibex/cs_registers_i/_1040_ ),
    .X(\i_ibex/cs_registers_i/mstatus_d [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/_2405_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/_1069_ ),
    .A(net624),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2406_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mstatus_q [3]),
    .A2(\i_ibex/cs_registers_i/mstatus_q [2]),
    .Y(\i_ibex/cs_registers_i/_1070_ ),
    .B1(\i_ibex/cs_registers_i/_1069_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2407_  (.A0(net943),
    .A1(\i_ibex/cs_registers_i/mstatus_q [1]),
    .S(net911),
    .X(\i_ibex/cs_registers_i/_1071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_2408_  (.A(\i_ibex/cs_registers_i/_1070_ ),
    .B_N(\i_ibex/cs_registers_i/_1071_ ),
    .Y(\i_ibex/cs_registers_i/mstatus_d [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout934 (.A(\i_ibex/cs_registers_i/csr_wdata_int [9]),
    .X(net934),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2411_  (.B(net482),
    .C(\i_ibex/cs_registers_i/_1040_ ),
    .A(\i_ibex/cs_registers_i/_1069_ ),
    .Y(\i_ibex/cs_registers_i/mstatus_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2412_  (.A0(\i_ibex/csr_mtval [31]),
    .A1(net422),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2413_  (.A0(\i_ibex/csr_mtval [30]),
    .A1(net963),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2415_  (.A0(\i_ibex/csr_mtval [21]),
    .A1(net961),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2416_  (.A0(\i_ibex/csr_mtval [20]),
    .A1(net426),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2417_  (.A0(\i_ibex/csr_mtval [19]),
    .A1(net947),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2418_  (.A0(\i_ibex/csr_mtval [18]),
    .A1(net945),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2419_  (.A0(\i_ibex/csr_mtval [17]),
    .A1(net943),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2420_  (.A0(\i_ibex/csr_mtval [16]),
    .A1(net941),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2421_  (.A0(\i_ibex/csr_mtval [15]),
    .A1(net960),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2422_  (.A(\i_ibex/csr_mtval [14]),
    .B(net482),
    .Y(\i_ibex/cs_registers_i/_1075_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2423_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0506_ ),
    .A2(net482),
    .Y(\i_ibex/cs_registers_i/mtval_d [14]),
    .B1(\i_ibex/cs_registers_i/_1075_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2424_  (.A0(\i_ibex/csr_mtval [13]),
    .A1(net958),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2425_  (.A0(\i_ibex/csr_mtval [12]),
    .A1(net939),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2426_  (.A0(\i_ibex/csr_mtval [29]),
    .A1(net420),
    .S(net478),
    .X(\i_ibex/cs_registers_i/mtval_d [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout932 (.A(\i_ibex/cs_registers_i/csr_wdata_int [8]),
    .X(net932),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2428_  (.A0(\i_ibex/csr_mtval [11]),
    .A1(net938),
    .S(net480),
    .X(\i_ibex/cs_registers_i/mtval_d [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2429_  (.A0(\i_ibex/csr_mtval [10]),
    .A1(net936),
    .S(net480),
    .X(\i_ibex/cs_registers_i/mtval_d [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2430_  (.A0(\i_ibex/csr_mtval [9]),
    .A1(net934),
    .S(net480),
    .X(\i_ibex/cs_registers_i/mtval_d [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2431_  (.A0(\i_ibex/csr_mtval [8]),
    .A1(net932),
    .S(net480),
    .X(\i_ibex/cs_registers_i/mtval_d [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2432_  (.A0(\i_ibex/csr_mtval [7]),
    .A1(net956),
    .S(net480),
    .X(\i_ibex/cs_registers_i/mtval_d [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2433_  (.A(\i_ibex/csr_mtval [6]),
    .B(net482),
    .Y(\i_ibex/cs_registers_i/_1077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2434_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0682_ ),
    .A2(net481),
    .Y(\i_ibex/cs_registers_i/mtval_d [6]),
    .B1(\i_ibex/cs_registers_i/_1077_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/_2435_  (.A(\i_ibex/csr_mtval [5]),
    .B(net481),
    .Y(\i_ibex/cs_registers_i/_1078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/_2436_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/_0195_ ),
    .A2(net481),
    .Y(\i_ibex/cs_registers_i/mtval_d [5]),
    .B1(\i_ibex/cs_registers_i/_1078_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2437_  (.A0(\i_ibex/csr_mtval [4]),
    .A1(net953),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2438_  (.A0(\i_ibex/csr_mtval [3]),
    .A1(net951),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2439_  (.A0(\i_ibex/csr_mtval [2]),
    .A1(net950),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2440_  (.A0(\i_ibex/csr_mtval [28]),
    .A1(net418),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2441_  (.A0(\i_ibex/csr_mtval [1]),
    .A1(net971),
    .S(net479),
    .X(\i_ibex/cs_registers_i/mtval_d [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2442_  (.A0(\i_ibex/csr_mtval [0]),
    .A1(net974),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2443_  (.A0(\i_ibex/csr_mtval [27]),
    .A1(net424),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2444_  (.A0(\i_ibex/csr_mtval [26]),
    .A1(net929),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2445_  (.A0(\i_ibex/csr_mtval [25]),
    .A1(net416),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2446_  (.A0(\i_ibex/csr_mtval [24]),
    .A1(net928),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2447_  (.A0(\i_ibex/csr_mtval [23]),
    .A1(net414),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2448_  (.A0(\i_ibex/csr_mtval [22]),
    .A1(net412),
    .S(net477),
    .X(\i_ibex/cs_registers_i/mtval_d [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/_2449_  (.B1(net481),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mtval_en ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/_0702_ ),
    .A2(\i_ibex/cs_registers_i/_1037_ ));
 sg13g2_buf_4 fanout931 (.X(net931),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2452_  (.A0(net422),
    .A1(net1771),
    .S(net1083),
    .X(\i_ibex/cs_registers_i/mtvec_d [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2453_  (.A0(net964),
    .A1(net1765),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2454_  (.A0(net962),
    .A1(net1775),
    .S(net1082),
    .X(\i_ibex/cs_registers_i/mtvec_d [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2455_  (.A0(net426),
    .A1(net1762),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2456_  (.A0(net947),
    .A1(net1778),
    .S(net1082),
    .X(\i_ibex/cs_registers_i/mtvec_d [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2457_  (.A0(net945),
    .A1(net1760),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2458_  (.A0(net944),
    .A1(net1773),
    .S(net1082),
    .X(\i_ibex/cs_registers_i/mtvec_d [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2459_  (.A0(net942),
    .A1(net1782),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2460_  (.A0(net960),
    .A1(net1780),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(net930),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2462_  (.A0(\i_ibex/cs_registers_i/csr_wdata_int [14]),
    .A1(net1783),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2463_  (.A0(net958),
    .A1(net1774),
    .S(net1084),
    .X(\i_ibex/cs_registers_i/mtvec_d [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2464_  (.A0(\i_ibex/cs_registers_i/csr_wdata_int [12]),
    .A1(net1764),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2465_  (.A0(net421),
    .A1(net1776),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2466_  (.A0(net938),
    .A1(net1763),
    .S(net1084),
    .X(\i_ibex/cs_registers_i/mtvec_d [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2467_  (.A0(net936),
    .A1(net1767),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2468_  (.A0(net934),
    .A1(net1761),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2469_  (.A0(net932),
    .A1(net1779),
    .S(net1084),
    .X(\i_ibex/cs_registers_i/mtvec_d [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2470_  (.A0(net418),
    .A1(net1777),
    .S(net1083),
    .X(\i_ibex/cs_registers_i/mtvec_d [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2471_  (.A0(net425),
    .A1(net1781),
    .S(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_d [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2472_  (.A0(net929),
    .A1(net1770),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2473_  (.A0(net416),
    .A1(net1759),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2474_  (.A0(net927),
    .A1(net1766),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2475_  (.A0(net414),
    .A1(net1768),
    .S(net1081),
    .X(\i_ibex/cs_registers_i/mtvec_d [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2476_  (.A0(net412),
    .A1(net1772),
    .S(net1083),
    .X(\i_ibex/cs_registers_i/mtvec_d [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/cs_registers_i/_2477_  (.A2(net926),
    .A1(net984),
    .B1(net1080),
    .X(\i_ibex/cs_registers_i/mtvec_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_2478_  (.A(\i_ibex/csr_save_cause ),
    .B_N(\i_ibex/cs_registers_i/_0000_ ),
    .Y(\i_ibex/cs_registers_i/_1082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2479_  (.A(\i_ibex/csr_restore_dret_id ),
    .B(net624),
    .C(\i_ibex/cs_registers_i/_1082_ ),
    .Y(\i_ibex/cs_registers_i/_1083_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_2480_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/mstatus_q [2]),
    .C1(\i_ibex/cs_registers_i/_1083_ ),
    .B1(net624),
    .A1(\i_ibex/csr_restore_dret_id ),
    .Y(\i_ibex/cs_registers_i/_0004_ ),
    .A2(\i_ibex/cs_registers_i/dcsr_q [0]));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/_2481_  (.A(\i_ibex/csr_save_cause ),
    .B_N(\i_ibex/cs_registers_i/_0001_ ),
    .Y(\i_ibex/cs_registers_i/_1084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/_2482_  (.A(\i_ibex/csr_restore_dret_id ),
    .B(net624),
    .C(\i_ibex/cs_registers_i/_1084_ ),
    .Y(\i_ibex/cs_registers_i/_1085_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/_2483_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net624),
    .C1(\i_ibex/cs_registers_i/_1085_ ),
    .B1(\i_ibex/cs_registers_i/mstatus_q [3]),
    .A1(\i_ibex/cs_registers_i/dcsr_q [1]),
    .Y(\i_ibex/cs_registers_i/_0005_ ),
    .A2(\i_ibex/csr_restore_dret_id ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2484_  (.A0(net785),
    .A1(\i_ibex/cs_registers_i/mstatus_q [3]),
    .S(\i_ibex/cs_registers_i/mstatus_q [1]),
    .X(\i_ibex/g_no_pmp.unused_priv_lvl_ls [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/_2485_  (.A0(net786),
    .A1(\i_ibex/cs_registers_i/mstatus_q [2]),
    .S(\i_ibex/cs_registers_i/mstatus_q [1]),
    .X(\i_ibex/g_no_pmp.unused_priv_lvl_ls [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2486_  (.Y(\i_ibex/cs_registers_i/_1086_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [5]),
    .B(\i_ibex/pc_if [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2487_  (.Y(\i_ibex/cs_registers_i/_1087_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [29]),
    .B(\i_ibex/pc_if [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2488_  (.Y(\i_ibex/cs_registers_i/_1088_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [10]),
    .B(\i_ibex/pc_if [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/_2489_  (.B(\i_ibex/cs_registers_i/_1087_ ),
    .C(\i_ibex/cs_registers_i/_1088_ ),
    .A(\i_ibex/cs_registers_i/_1086_ ),
    .Y(\i_ibex/cs_registers_i/_1089_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2490_  (.Y(\i_ibex/cs_registers_i/_1090_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [19]),
    .B(\i_ibex/pc_if [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2491_  (.Y(\i_ibex/cs_registers_i/_1091_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [1]),
    .B(net1478),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2492_  (.Y(\i_ibex/cs_registers_i/_1092_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [18]),
    .B(\i_ibex/pc_if [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2493_  (.Y(\i_ibex/cs_registers_i/_1093_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [6]),
    .B(\i_ibex/pc_if [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2494_  (.B(\i_ibex/cs_registers_i/_1091_ ),
    .C(\i_ibex/cs_registers_i/_1092_ ),
    .A(\i_ibex/cs_registers_i/_1090_ ),
    .Y(\i_ibex/cs_registers_i/_1094_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1093_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2495_  (.Y(\i_ibex/cs_registers_i/_1095_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [13]),
    .B(\i_ibex/pc_if [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2496_  (.Y(\i_ibex/cs_registers_i/_1096_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [28]),
    .B(\i_ibex/pc_if [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2497_  (.Y(\i_ibex/cs_registers_i/_1097_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [23]),
    .B(\i_ibex/pc_if [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2498_  (.Y(\i_ibex/cs_registers_i/_1098_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [31]),
    .B(\i_ibex/pc_if [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2499_  (.B(\i_ibex/cs_registers_i/_1096_ ),
    .C(\i_ibex/cs_registers_i/_1097_ ),
    .A(\i_ibex/cs_registers_i/_1095_ ),
    .Y(\i_ibex/cs_registers_i/_1099_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1098_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2500_  (.Y(\i_ibex/cs_registers_i/_1100_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [11]),
    .B(\i_ibex/pc_if [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/_2501_  (.B(\i_ibex/pc_if [2]),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [2]),
    .X(\i_ibex/cs_registers_i/_1101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/_2502_  (.B(\i_ibex/pc_if [15]),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [15]),
    .X(\i_ibex/cs_registers_i/_1102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/_2503_  (.B(\i_ibex/pc_if [24]),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [24]),
    .X(\i_ibex/cs_registers_i/_1103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/_2504_  (.B(\i_ibex/pc_if [12]),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [12]),
    .X(\i_ibex/cs_registers_i/_1104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_2505_  (.A(\i_ibex/cs_registers_i/_1101_ ),
    .B(\i_ibex/cs_registers_i/_1102_ ),
    .C(\i_ibex/cs_registers_i/_1103_ ),
    .D(\i_ibex/cs_registers_i/_1104_ ),
    .Y(\i_ibex/cs_registers_i/_1105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2506_  (.Y(\i_ibex/cs_registers_i/_1106_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [27]),
    .B(\i_ibex/pc_if [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2507_  (.Y(\i_ibex/cs_registers_i/_1107_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [21]),
    .B(\i_ibex/pc_if [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2508_  (.Y(\i_ibex/cs_registers_i/_1108_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [25]),
    .B(\i_ibex/pc_if [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2509_  (.Y(\i_ibex/cs_registers_i/_1109_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [17]),
    .B(\i_ibex/pc_if [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2510_  (.B(\i_ibex/cs_registers_i/_1107_ ),
    .C(\i_ibex/cs_registers_i/_1108_ ),
    .A(\i_ibex/cs_registers_i/_1106_ ),
    .Y(\i_ibex/cs_registers_i/_1110_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1109_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2511_  (.Y(\i_ibex/cs_registers_i/_1111_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [0]),
    .B(net379),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2512_  (.Y(\i_ibex/cs_registers_i/_1112_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [16]),
    .B(\i_ibex/pc_if [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2513_  (.Y(\i_ibex/cs_registers_i/_1113_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [14]),
    .B(\i_ibex/pc_if [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2514_  (.Y(\i_ibex/cs_registers_i/_1114_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [9]),
    .B(\i_ibex/pc_if [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2515_  (.B(\i_ibex/cs_registers_i/_1112_ ),
    .C(\i_ibex/cs_registers_i/_1113_ ),
    .A(\i_ibex/cs_registers_i/_1111_ ),
    .Y(\i_ibex/cs_registers_i/_1115_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1114_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2516_  (.Y(\i_ibex/cs_registers_i/_1116_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [26]),
    .B(\i_ibex/pc_if [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2517_  (.Y(\i_ibex/cs_registers_i/_1117_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [8]),
    .B(\i_ibex/pc_if [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2518_  (.Y(\i_ibex/cs_registers_i/_1118_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [3]),
    .B(\i_ibex/pc_if [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2519_  (.Y(\i_ibex/cs_registers_i/_1119_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [20]),
    .B(\i_ibex/pc_if [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2520_  (.B(\i_ibex/cs_registers_i/_1117_ ),
    .C(\i_ibex/cs_registers_i/_1118_ ),
    .A(\i_ibex/cs_registers_i/_1116_ ),
    .Y(\i_ibex/cs_registers_i/_1120_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1119_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2521_  (.Y(\i_ibex/cs_registers_i/_1121_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [22]),
    .B(\i_ibex/pc_if [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2522_  (.Y(\i_ibex/cs_registers_i/_1122_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [7]),
    .B(\i_ibex/pc_if [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2523_  (.Y(\i_ibex/cs_registers_i/_1123_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [30]),
    .B(\i_ibex/pc_if [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/_2524_  (.Y(\i_ibex/cs_registers_i/_1124_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [4]),
    .B(\i_ibex/pc_if [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2525_  (.B(\i_ibex/cs_registers_i/_1122_ ),
    .C(\i_ibex/cs_registers_i/_1123_ ),
    .A(\i_ibex/cs_registers_i/_1121_ ),
    .Y(\i_ibex/cs_registers_i/_1125_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1124_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/_2526_  (.A(\i_ibex/cs_registers_i/_1110_ ),
    .B(\i_ibex/cs_registers_i/_1115_ ),
    .C(\i_ibex/cs_registers_i/_1120_ ),
    .D(\i_ibex/cs_registers_i/_1125_ ),
    .Y(\i_ibex/cs_registers_i/_1126_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/_2527_  (.B(\i_ibex/cs_registers_i/_1100_ ),
    .C(\i_ibex/cs_registers_i/_1105_ ),
    .A(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_control ),
    .Y(\i_ibex/cs_registers_i/_1127_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1126_ ));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/_2528_  (.A(\i_ibex/cs_registers_i/_1089_ ),
    .B(\i_ibex/cs_registers_i/_1094_ ),
    .C(\i_ibex/cs_registers_i/_1099_ ),
    .Y(\i_ibex/trigger_match ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/_1127_ ));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(net474),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1474__72  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net72));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/_3_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_control ),
    .A1(net949),
    .S(\i_ibex/cs_registers_i/gen_trigger_regs.tmatch_control_we ),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/_0_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1458__71  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net71));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/rd_data_o_reg  (.CLK(clknet_leaf_45_clk_i_regs),
    .RESET_B(net1606),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/_0_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr/_1_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_control ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(net928),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_071_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [0]),
    .A1(net973),
    .S(net886),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_072_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [10]),
    .A1(net936),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_073_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [11]),
    .A1(net937),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_074_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [12]),
    .A1(net939),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_075_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [13]),
    .A1(net958),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_076_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [14]),
    .A1(net940),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_077_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [15]),
    .A1(net959),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_078_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [16]),
    .A1(net941),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_079_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [17]),
    .A1(net943),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_080_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [18]),
    .A1(net945),
    .S(net888),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(\i_ibex/cs_registers_i/_0864_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_082_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [19]),
    .A1(net947),
    .S(net888),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_083_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [1]),
    .A1(net972),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_084_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [20]),
    .A1(net426),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_085_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [21]),
    .A1(net961),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_086_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [22]),
    .A1(net412),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_087_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [23]),
    .A1(net414),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_088_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [24]),
    .A1(net927),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_089_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [25]),
    .A1(net416),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_090_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [26]),
    .A1(net929),
    .S(net887),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_091_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [27]),
    .A1(net424),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(\i_ibex/cs_registers_i/depc_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_093_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [28]),
    .A1(net418),
    .S(net888),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_094_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [29]),
    .A1(net420),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_095_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [2]),
    .A1(net950),
    .S(net886),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_096_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [30]),
    .A1(net963),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_097_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [31]),
    .A1(net422),
    .S(net888),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_098_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [3]),
    .A1(net951),
    .S(net886),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_099_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [4]),
    .A1(net954),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_100_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [5]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_101_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [6]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_102_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [7]),
    .A1(net956),
    .S(net886),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_103_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [8]),
    .A1(net931),
    .S(net889),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_104_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [9]),
    .A1(net933),
    .S(net885),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1457__70  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net70));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[0]_reg  (.RESET_B(net1605),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_000_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [0]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_067_ ),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_45_clk_i_regs),
    .RESET_B(net1605),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_001_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_46_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_065_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[12]_reg  (.RESET_B(net1599),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_003_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [12]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_064_ ),
    .CLK(clknet_leaf_51_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[13]_reg  (.RESET_B(net1636),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_004_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [13]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_063_ ),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_46_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_47_clk_i_regs),
    .RESET_B(net1636),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_24_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[1]_reg  (.RESET_B(net1538),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_011_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [1]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_056_ ),
    .CLK(clknet_leaf_77_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1590),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_24_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[22]_reg  (.RESET_B(net1617),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_014_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [22]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_053_ ),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[23]_reg  (.RESET_B(net1617),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_015_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [23]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_052_ ),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_25_clk_i_regs),
    .RESET_B(net1617),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[25]_reg  (.RESET_B(net1617),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_017_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [25]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_050_ ),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[26]_reg  (.RESET_B(net1619),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_018_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [26]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_049_ ),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_21_clk_i_regs),
    .RESET_B(net1590),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[28]_reg  (.RESET_B(net1631),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_020_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [28]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_047_ ),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[29]_reg  (.RESET_B(net1595),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_021_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [29]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_046_ ),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_79_clk_i_regs),
    .RESET_B(net1610),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_045_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[30]_reg  (.RESET_B(net1621),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_023_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [30]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_044_ ),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1630),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_043_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_79_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[4]_reg  (.RESET_B(net1538),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_026_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [4]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_041_ ),
    .CLK(clknet_leaf_77_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[5]_reg  (.RESET_B(net1531),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_027_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [5]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_040_ ),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[6]_reg  (.RESET_B(net1529),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_028_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [6]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_039_ ),
    .CLK(clknet_leaf_60_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[7]_reg  (.RESET_B(net1531),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_029_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [7]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_038_ ),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[8]_reg  (.RESET_B(net1604),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_030_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [8]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_037_ ),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/rd_data_o[9]_reg  (.RESET_B(net1600),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_031_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.selected_tmatch_value [9]),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr/_036_ ),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_3_  (.A0(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_q ),
    .A1(net46),
    .S(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_we ),
    .X(\i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_0_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1449__69  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net69));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/rd_data_o_reg  (.CLK(clknet_leaf_45_clk_i_regs),
    .RESET_B(net1605),
    .D(\i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_0_ ),
    .Q_N(\i_ibex/cs_registers_i/gen_trigger_regs.u_tselect_csr/_1_ ),
    .Q(\i_ibex/cs_registers_i/gen_trigger_regs.tselect_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcountinhibit[0]_reg  (.RESET_B(net1534),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/_0002_ ),
    .Q(\i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y [192]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .CLK(clknet_leaf_65_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcountinhibit[2]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1539),
    .D(\i_ibex/cs_registers_i/_0003_ ),
    .Q_N(\i_ibex/cs_registers_i/instr_ret_i_$_AND__A_B ),
    .Q(\i_ibex/cs_registers_i/irq_timer_i_$_AND__A_Y_$_NOT__Y_1_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y [194]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(net925),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout923 (.A(net925),
    .X(net923),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(net923),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout921 (.A(net925),
    .X(net921),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net925),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout919 (.A(\i_ibex/cs_registers_i/mhpmcounter_we [0]),
    .X(net919),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout918 (.A(net919),
    .X(net918),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/mcycle_counter_i/_408_  (.A(net919),
    .B_N(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_409_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_072_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_071_ ),
    .B2(\i_ibex/cs_registers_i/mcycle_counter_i/counter_upd [0]),
    .A2(net915),
    .A1(net973),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout917 (.X(net917),
    .A(net918),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout916 (.X(net916),
    .A(net917),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_412_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .B(net915),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_075_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_413_  (.B1(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_076_ ),
    .VSS(VSS),
    .A1(net401),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_075_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_414_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_076_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_000_ ),
    .VSS(VSS),
    .A1(net400),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_072_ ));
 sg13g2_buf_2 fanout915 (.A(net919),
    .X(net915),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_416_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1986]),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_078_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [1985]));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_417_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1989]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1988]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1990]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [1987]));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/mcycle_counter_i/_418_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_078_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_079_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/mcycle_counter_i/_419_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1991]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_420_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_082_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1993]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [1992]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_421_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_083_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_082_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ));
 sg13g2_buf_2 fanout914 (.A(net919),
    .X(net914),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_423_  (.A(net403),
    .B(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_082_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_085_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_424_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_083_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_086_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_085_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_425_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_087_ ),
    .A(net914),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_426_  (.A(net406),
    .B(net863),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout913 (.A(net914),
    .X(net913),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_428_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_090_ ),
    .B1(net850),
    .B2(net935),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .A1(net405),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_429_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_090_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_001_ ),
    .VSS(VSS),
    .A1(net914),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_086_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_430_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_091_ ),
    .A(net405),
    .VSS(VSS));
 sg13g2_buf_2 fanout912 (.A(net914),
    .X(net912),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/cs_registers_i/mcycle_counter_i/_432_  (.B(net397),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_093_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/cs_registers_i/mcycle_counter_i/_083_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_433_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1995]),
    .B(net850),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_094_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_434_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_095_ ),
    .A(net395),
    .B(net918),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout911 (.A(\i_ibex/cs_registers_i/_1040_ ),
    .X(net911),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_436_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1993]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1995]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_097_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [1992]));
 sg13g2_or4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_437_  (.A(net406),
    .B(net915),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_097_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_438_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_098_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_099_ ),
    .VSS(VSS),
    .A1(net937),
    .A2(net862));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_439_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_093_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_094_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_002_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_099_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_440_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_100_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_097_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_441_  (.A(net403),
    .B(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_097_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_442_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_100_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_102_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_101_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_443_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_103_ ),
    .B1(net850),
    .B2(net939),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .A1(net405),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_444_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_103_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_003_ ),
    .VSS(VSS),
    .A1(net915),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_102_ ));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_445_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1997]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_446_  (.A0(net957),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1997]),
    .S(net862),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_447_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_104_ ),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_105_ ),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_098_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_448_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_106_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1997]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_449_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_107_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1998]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_450_  (.A0(net940),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1998]),
    .S(net862),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_451_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_107_ ),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_108_ ),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_098_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_452_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1997]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1998]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_109_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [1991]));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_453_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_078_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_079_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_097_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_110_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_109_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_454_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .B(net918),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_455_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_112_ ),
    .B1(net695),
    .B2(\i_ibex/cs_registers_i/mcycle_counter_i/_111_ ),
    .A2(net918),
    .A1(net959),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_456_  (.B1(net395),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_113_ ),
    .VSS(VSS),
    .A1(net918),
    .A2(net695));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_457_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_114_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_458_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_114_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_006_ ),
    .VSS(VSS),
    .A1(net400),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_112_ ));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_459_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .C(net863),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2000]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_115_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net695));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_460_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_115_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_116_ ),
    .VSS(VSS),
    .A1(net942),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_087_ ));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/mcycle_counter_i/_461_  (.A2(net695),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .B1(net916),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_117_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_462_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net396),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_117_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_118_ ),
    .B1(\i_ibex/cs_registers_i/mhpmcounter [2000]));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_463_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net396),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_116_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_007_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_118_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_464_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2001]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_115_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_465_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net943),
    .A2(net916),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_120_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_119_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_466_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .C(net695),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2000]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_467_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_087_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_121_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_122_ ),
    .B1(net402));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/mcycle_counter_i/_468_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_123_ ),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2001]),
    .A_N(\i_ibex/cs_registers_i/mcycle_counter_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_469_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_123_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_008_ ),
    .VSS(VSS),
    .A1(net400),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_120_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_470_  (.A(net406),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2002]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_471_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2000]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2001]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_125_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net695));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_472_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_124_ ),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2002]),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_125_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_126_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_473_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_127_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_126_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_474_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_128_ ),
    .B1(net849),
    .B2(net946),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2002]),
    .A1(net405),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_475_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_128_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_009_ ),
    .VSS(VSS),
    .A1(net917),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_127_ ));
 sg13g2_and4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_476_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2002]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2001]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2000]),
    .D(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/mcycle_counter_i/_477_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .A(net695),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_478_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .B(net916),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_479_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net948),
    .A2(net917),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_132_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_131_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_480_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net695),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_129_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_133_ ),
    .B1(net916));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_481_  (.B1(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_134_ ),
    .VSS(VSS),
    .A1(net401),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_133_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_482_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_134_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_010_ ),
    .VSS(VSS),
    .A1(net400),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_132_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_483_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_135_ ),
    .A(net971),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_484_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1985]),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_485_  (.A(net912),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_136_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_486_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_135_ ),
    .A2(net913),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_138_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_137_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_487_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_139_ ),
    .B1(net915));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_488_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_140_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1985]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_489_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_140_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_141_ ),
    .VSS(VSS),
    .A1(net402),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_139_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_490_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_141_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_142_ ),
    .VSS(VSS),
    .A1(net400),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_138_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_491_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_011_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_142_ ),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_492_  (.A(net426),
    .B(net850),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_143_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_493_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2004]),
    .A2(net862),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_144_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_143_ ));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/mcycle_counter_i/_494_  (.A(net405),
    .B(net916),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_495_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_097_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_109_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_146_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_496_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_145_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_146_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_080_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_129_ ));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_497_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2004]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_148_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_498_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_148_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_149_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_499_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_144_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_012_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_149_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_500_  (.A(net961),
    .B(net850),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_501_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2005]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_151_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_150_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_502_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_152_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2004]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_503_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_153_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2005]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_152_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_504_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_153_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_505_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_151_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_013_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_154_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_506_  (.A(net412),
    .B(net850),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_507_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2006]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_156_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_155_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_508_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2004]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2005]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_509_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_158_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2006]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_510_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_158_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_511_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_156_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_014_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_159_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_512_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_160_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2007]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2006]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_513_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_157_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_514_  (.A0(net414),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2007]),
    .S(net861),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_162_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_515_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_162_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_161_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_516_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_160_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_161_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_015_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_163_ ));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(\i_ibex/cs_registers_i/_0866_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_518_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_165_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2007]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2006]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_519_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_157_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_165_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_166_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_520_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_129_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_166_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_110_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_521_  (.A(net402),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_167_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_522_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_167_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_169_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_168_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_523_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_170_ ),
    .B1(net849),
    .B2(net928),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .A1(net405),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_524_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_170_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_016_ ),
    .VSS(VSS),
    .A1(net916),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_169_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_525_  (.A(net416),
    .B(net849),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_171_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_526_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_172_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_171_ ));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/mcycle_counter_i/_527_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_173_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_166_ ),
    .A_N(\i_ibex/cs_registers_i/mcycle_counter_i/_147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_528_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_174_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_529_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_174_ ),
    .B(net848),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_530_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_172_ ),
    .A2(net848),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_017_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_175_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_531_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_176_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_532_  (.B1(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_177_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_167_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_176_ ));
 sg13g2_or4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_533_  (.A(net405),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_167_ ),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_176_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_534_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_177_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_178_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_179_ ),
    .B1(net916));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_535_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_180_ ),
    .B1(net849),
    .B2(net930),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .A1(net405),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/mcycle_counter_i/_536_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_018_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_180_ ),
    .A_N(\i_ibex/cs_registers_i/mcycle_counter_i/_179_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_537_  (.A(net424),
    .B(net849),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_181_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_538_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2011]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_182_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_181_ ));
 sg13g2_and3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_539_  (.X(\i_ibex/cs_registers_i/mcycle_counter_i/_183_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_540_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_183_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2011]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_541_  (.A(net848),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_184_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_542_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net848),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_182_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_019_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_185_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_543_  (.A(net418),
    .B(net849),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_186_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_544_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2012]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_187_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_186_ ));
 sg13g2_and4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_545_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2011]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .D(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_546_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_188_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2012]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_547_  (.A(net848),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_189_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_548_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net848),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_187_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_020_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_190_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_549_  (.A(net420),
    .B(net849),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_191_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_550_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2013]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_192_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_191_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_551_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2011]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_183_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2012]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_552_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_194_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2013]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_553_  (.A(net848),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_194_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_195_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_554_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net848),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_192_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_021_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_195_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_555_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_196_ ),
    .A(net949),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_556_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_197_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_137_ ),
    .B2(\i_ibex/cs_registers_i/mhpmcounter [1986]),
    .A2(net913),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_557_  (.A(net406),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_197_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_558_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net863),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_136_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_199_ ),
    .B1(net402));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_559_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1986]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_199_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_560_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_198_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_200_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_561_  (.A(net963),
    .B(net849),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_201_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_562_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [2014]),
    .A2(net861),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_202_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_201_ ));
 sg13g2_and3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_563_  (.X(\i_ibex/cs_registers_i/mcycle_counter_i/_203_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2013]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2012]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_564_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_203_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2014]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_565_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_173_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_204_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_566_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_173_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_202_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_023_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_205_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_567_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_206_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2015]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_568_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_207_ ),
    .A(net395),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_206_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_569_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_208_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2014]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_570_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_157_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_165_ ),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_208_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_571_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_206_ ),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_207_ ),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_209_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_210_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_572_  (.X(\i_ibex/cs_registers_i/mcycle_counter_i/_211_ ),
    .A(net395),
    .B(net422),
    .C(net917),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_573_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net406),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2015]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_212_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_211_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_574_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_212_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_024_ ),
    .VSS(VSS),
    .A1(net917),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_210_ ));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_575_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_206_ ),
    .B(net916),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_167_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_213_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_208_ ));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_576_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_213_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2016]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_214_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_577_  (.A0(net973),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_214_ ),
    .S(net397),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_578_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_215_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2017]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2016]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_579_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_145_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_166_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2014]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_216_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_203_ ));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/mcycle_counter_i/_580_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_206_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .C(net1515),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_581_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2017]),
    .A1(net971),
    .S(net401),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_218_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_582_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_218_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_219_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_583_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_215_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_026_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_219_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_584_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2018]),
    .A1(net949),
    .S(net401),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_220_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_585_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_221_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2017]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2016]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_586_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_222_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2018]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_221_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_587_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_220_ ),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_222_ ),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_588_  (.X(\i_ibex/cs_registers_i/mcycle_counter_i/_223_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2018]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2017]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2016]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_589_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_224_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_590_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2019]),
    .A1(net952),
    .S(net402),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_591_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_028_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_224_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_592_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2020]),
    .A1(net953),
    .S(net401),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_226_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_593_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_227_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2019]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_594_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_228_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2020]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_595_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_226_ ),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_228_ ),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_596_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2019]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2020]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_229_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_223_ ));
 sg13g2_buf_2 fanout909 (.A(net910),
    .X(net909),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_598_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2021]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .S(net404),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_599_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_030_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_229_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_600_  (.X(\i_ibex/cs_registers_i/mcycle_counter_i/_232_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2021]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2020]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2019]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_601_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_223_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_232_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_602_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_234_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_603_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2022]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .S(net404),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_235_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_604_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_031_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_234_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_235_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_605_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_217_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_233_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2022]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_236_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_606_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2023]),
    .A1(net955),
    .S(net404),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_607_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_032_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_236_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_608_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i_counter_inc_i ),
    .B(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1986]),
    .D(\i_ibex/cs_registers_i/mhpmcounter [1985]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_238_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_609_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .B(net912),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_239_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_610_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_240_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_238_ ),
    .B2(\i_ibex/cs_registers_i/mcycle_counter_i/_239_ ),
    .A2(net912),
    .A1(net952),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_611_  (.B1(net395),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_241_ ),
    .VSS(VSS),
    .A1(net913),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_238_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_612_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_242_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_241_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_613_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_242_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_033_ ),
    .VSS(VSS),
    .A1(net400),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_240_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_614_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2023]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2015]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_243_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_615_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_223_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_232_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2022]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_244_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_243_ ));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/mcycle_counter_i/_616_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .B(net1515),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_244_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_245_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_617_  (.A(net398),
    .B(net931),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_618_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net396),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2024]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_247_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_246_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_619_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_034_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_245_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_620_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_248_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2024]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_245_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_621_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2025]),
    .A1(net933),
    .S(net404),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_249_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_622_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_035_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_248_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_249_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_623_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2024]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_245_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2025]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_250_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_624_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2026]),
    .A1(net935),
    .S(net403),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_625_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_036_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_250_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_626_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2025]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2024]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2026]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_252_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_245_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_627_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2027]),
    .A1(net937),
    .S(net403),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_628_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_037_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_252_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_629_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2026]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2025]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2027]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [2024]));
 sg13g2_or2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_630_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_255_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_254_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_244_ ));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/mcycle_counter_i/_631_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .B(net1515),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_255_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_256_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_632_  (.A(net398),
    .B(net939),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_257_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_633_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net396),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2028]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_258_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_257_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_634_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_038_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_256_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_635_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_259_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2028]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_256_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_636_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2029]),
    .A1(net957),
    .S(net403),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_637_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_039_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_259_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_638_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2028]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_256_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2029]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_639_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2030]),
    .A1(net940),
    .S(net403),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_640_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_040_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_261_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_641_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2029]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2028]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2030]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_263_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_256_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_642_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2031]),
    .A1(net959),
    .S(net403),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_643_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_041_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_263_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_644_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2030]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2029]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2031]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_265_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [2028]));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_645_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .B(net1515),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_255_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_265_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_646_  (.A(net398),
    .B(net942),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_267_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_647_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net396),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2032]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_268_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_267_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_648_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_042_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_266_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_649_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_269_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2032]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_650_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2033]),
    .A1(net943),
    .S(net403),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_270_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_651_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_043_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_269_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_270_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_652_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_238_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1988]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_271_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_653_  (.A0(net953),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_271_ ),
    .S(net863),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_272_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_654_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_238_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_273_ ),
    .B1(net912));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_655_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_274_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1988]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_656_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_274_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_275_ ),
    .VSS(VSS),
    .A1(net402),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_273_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_657_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_275_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_276_ ),
    .VSS(VSS),
    .A1(net401),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_272_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_658_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_044_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_276_ ),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_659_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2032]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_266_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2033]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_277_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_660_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2034]),
    .A1(net946),
    .S(net399),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_661_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_045_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_277_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_662_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2035]),
    .A1(net948),
    .S(net399),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_279_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_663_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2033]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2032]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2034]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_280_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_266_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_664_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_046_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_279_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_280_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_665_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2034]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2033]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2035]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_281_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mhpmcounter [2032]));
 sg13g2_or4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_666_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_244_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_254_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_265_ ),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_281_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_282_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/mcycle_counter_i/_667_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_216_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_282_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_283_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_668_  (.A(net398),
    .B(net426),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_284_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_669_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net395),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_285_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_284_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_670_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_047_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_283_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_285_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_671_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2037]),
    .A1(net961),
    .S(net399),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_286_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_672_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_287_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_283_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_673_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_048_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_286_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_287_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_674_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2038]),
    .A1(net412),
    .S(net399),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_288_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_675_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_283_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2037]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_289_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_676_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_049_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_288_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_289_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_677_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2039]),
    .A1(net414),
    .S(net399),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_290_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_678_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2038]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2037]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_291_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_283_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_679_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_050_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_290_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_291_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_680_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2040]),
    .A1(net928),
    .S(net399),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_292_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_681_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2037]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [2039]),
    .D(\i_ibex/cs_registers_i/mhpmcounter [2038]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_682_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_294_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_283_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_683_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_051_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_292_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_294_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_684_  (.A(net398),
    .B(net416),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_685_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net395),
    .A2(\i_ibex/cs_registers_i/mhpmcounter [2041]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_296_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_295_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_686_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_297_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2040]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/mcycle_counter_i/_687_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_130_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_216_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_282_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_297_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_688_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_052_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_296_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_689_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2042]),
    .A1(net930),
    .S(net398),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_299_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_690_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_300_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2041]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_691_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_053_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_299_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_692_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2043]),
    .A1(net424),
    .S(net398),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_301_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_693_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2042]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2041]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_694_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_303_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_695_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_054_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_301_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_696_  (.B(\i_ibex/cs_registers_i/mhpmcounter [1988]),
    .C(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1989]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_304_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_238_ ));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/mcycle_counter_i/_697_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_305_ ),
    .B(net912),
    .A_N(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_698_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_305_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_306_ ),
    .VSS(VSS),
    .A1(net912),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_304_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_699_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net863),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_271_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_307_ ),
    .B1(net402));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_700_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1989]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_307_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_308_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_701_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net396),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_306_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_055_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_308_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_702_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2044]),
    .A1(net418),
    .S(net401),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_309_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_703_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_302_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2043]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_704_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_056_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_309_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_705_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2045]),
    .A1(net420),
    .S(net400),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_311_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_706_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2043]),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2044]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_312_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_302_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_707_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_057_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_311_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_708_  (.A(\i_ibex/cs_registers_i/mhpmcounter [2045]),
    .B(\i_ibex/cs_registers_i/mhpmcounter [2044]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_709_  (.B(\i_ibex/cs_registers_i/mcycle_counter_i/_298_ ),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_302_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2043]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_314_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_313_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_710_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2046]),
    .A1(net963),
    .S(net398),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_711_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_058_ ),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_314_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_712_  (.B(\i_ibex/cs_registers_i/mhpmcounter [2046]),
    .A(\i_ibex/cs_registers_i/mhpmcounter [2047]),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_316_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_713_  (.A0(\i_ibex/cs_registers_i/mhpmcounter [2047]),
    .A1(net422),
    .S(net400),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_317_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_714_  (.A0(\i_ibex/cs_registers_i/mcycle_counter_i/_316_ ),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_317_ ),
    .S(\i_ibex/cs_registers_i/mcycle_counter_i/_314_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_715_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_318_ ),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_716_  (.A(net912),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_304_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_717_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_320_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_319_ ),
    .B2(\i_ibex/cs_registers_i/mhpmcounter [1990]),
    .A2(net912),
    .A1(\i_ibex/cs_registers_i/mcycle_counter_i/_318_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_718_  (.A(net406),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_320_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_719_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net863),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_304_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_322_ ),
    .B1(net402));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_720_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1990]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_322_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_721_  (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_321_ ),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_323_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_060_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_722_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1991]),
    .B(net915),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_324_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_723_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_325_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_080_ ),
    .B2(\i_ibex/cs_registers_i/mcycle_counter_i/_324_ ),
    .A2(net915),
    .A1(net955),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_724_  (.B1(net396),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_326_ ),
    .VSS(VSS),
    .A1(net915),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_080_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_725_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_327_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1991]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_326_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_726_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_327_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_061_ ),
    .VSS(VSS),
    .A1(net399),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_325_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/mcycle_counter_i/_727_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1991]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_080_ ),
    .X(\i_ibex/cs_registers_i/mcycle_counter_i/_328_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/mcycle_counter_i/_728_  (.B(net863),
    .C(\i_ibex/cs_registers_i/mcycle_counter_i/_328_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1992]),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_729_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_329_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_330_ ),
    .VSS(VSS),
    .A1(net931),
    .A2(net863));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_730_  (.B1(net396),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_331_ ),
    .VSS(VSS),
    .A1(net914),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_328_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/mcycle_counter_i/_731_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_332_ ),
    .A(\i_ibex/cs_registers_i/mhpmcounter [1992]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_732_  (.Y(\i_ibex/cs_registers_i/mcycle_counter_i/_062_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_331_ ),
    .B2(\i_ibex/cs_registers_i/mcycle_counter_i/_332_ ),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_330_ ),
    .A1(net395),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/mcycle_counter_i/_733_  (.A(\i_ibex/cs_registers_i/mhpmcounter [1993]),
    .B(\i_ibex/cs_registers_i/mcycle_counter_i/_332_ ),
    .C(net914),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_081_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_333_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_734_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net933),
    .A2(net913),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_334_ ),
    .B1(\i_ibex/cs_registers_i/mcycle_counter_i/_333_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/mcycle_counter_i/_735_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mhpmcounter [1992]),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_328_ ),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_335_ ),
    .B1(net913));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_736_  (.B1(\i_ibex/cs_registers_i/mhpmcounter [1993]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_336_ ),
    .VSS(VSS),
    .A1(net401),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_335_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/mcycle_counter_i/_737_  (.B1(\i_ibex/cs_registers_i/mcycle_counter_i/_336_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/mcycle_counter_i/_063_ ),
    .VSS(VSS),
    .A1(net399),
    .A2(\i_ibex/cs_registers_i/mcycle_counter_i/_334_ ));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1448__68  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net68));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[0]_reg  (.RESET_B(net1528),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_000_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1984]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/counter_upd [0]),
    .CLK(clknet_leaf_59_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[10]_reg  (.RESET_B(net1530),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_001_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1994]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_399_ ),
    .CLK(clknet_leaf_56_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[11]_reg  (.CLK(clknet_leaf_56_clk_i_regs),
    .RESET_B(net1530),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_398_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1995]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[12]_reg  (.RESET_B(net1529),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_003_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1996]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_397_ ),
    .CLK(clknet_leaf_56_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[13]_reg  (.RESET_B(net1530),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_004_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1997]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_396_ ),
    .CLK(clknet_leaf_51_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[14]_reg  (.CLK(clknet_leaf_51_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_395_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1998]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[15]_reg  (.RESET_B(net1589),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_006_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1999]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_394_ ),
    .CLK(clknet_leaf_53_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[16]_reg  (.RESET_B(net1590),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_007_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2000]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_393_ ),
    .CLK(clknet_leaf_53_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[17]_reg  (.CLK(clknet_leaf_53_clk_i_regs),
    .RESET_B(net1590),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_392_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2001]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[18]_reg  (.CLK(clknet_leaf_17_clk_i_regs),
    .RESET_B(net1590),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_391_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2002]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[19]_reg  (.RESET_B(net1590),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_010_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2003]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_390_ ),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[1]_reg  (.CLK(clknet_leaf_65_clk_i_regs),
    .RESET_B(net1534),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_389_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1985]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[20]_reg  (.RESET_B(net1587),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_012_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2004]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_388_ ),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[21]_reg  (.CLK(clknet_leaf_18_clk_i_regs),
    .RESET_B(net1587),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_387_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2005]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[22]_reg  (.RESET_B(net1587),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_014_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2006]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_386_ ),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[23]_reg  (.CLK(clknet_leaf_18_clk_i_regs),
    .RESET_B(net1597),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_385_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2007]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[24]_reg  (.RESET_B(net1587),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_016_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2008]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_384_ ),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[25]_reg  (.RESET_B(net1585),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_017_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2009]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_383_ ),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[26]_reg  (.RESET_B(net1585),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_018_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2010]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_382_ ),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[27]_reg  (.RESET_B(net1585),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_019_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2011]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_381_ ),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[28]_reg  (.RESET_B(net1585),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_020_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2012]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_380_ ),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[29]_reg  (.CLK(clknet_leaf_15_clk_i_regs),
    .RESET_B(net1586),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_379_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2013]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[2]_reg  (.RESET_B(net1534),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_022_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1986]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_378_ ),
    .CLK(clknet_leaf_65_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[30]_reg  (.RESET_B(net1586),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_023_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2014]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_377_ ),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[31]_reg  (.RESET_B(net1590),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_024_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2015]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_376_ ),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[32]_reg  (.RESET_B(net1530),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_025_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2016]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_375_ ),
    .CLK(clknet_leaf_55_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[33]_reg  (.RESET_B(net1540),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_026_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2017]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_374_ ),
    .CLK(clknet_leaf_69_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[34]_reg  (.RESET_B(net1544),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_027_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2018]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_373_ ),
    .CLK(clknet_leaf_69_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[35]_reg  (.RESET_B(net1540),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_028_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2019]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_372_ ),
    .CLK(clknet_leaf_67_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[36]_reg  (.RESET_B(net1540),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_029_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2020]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_371_ ),
    .CLK(clknet_leaf_69_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[37]_reg  (.CLK(clknet_leaf_67_clk_i_regs),
    .RESET_B(net1535),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_370_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2021]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[38]_reg  (.CLK(clknet_leaf_67_clk_i_regs),
    .RESET_B(net1535),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_369_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2022]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[39]_reg  (.CLK(clknet_leaf_67_clk_i_regs),
    .RESET_B(net1535),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_032_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_368_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2023]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[3]_reg  (.RESET_B(net1534),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_033_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1987]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_367_ ),
    .CLK(clknet_leaf_65_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[40]_reg  (.RESET_B(net1601),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_034_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2024]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_366_ ),
    .CLK(clknet_leaf_57_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[41]_reg  (.RESET_B(net1528),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_035_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2025]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_365_ ),
    .CLK(clknet_leaf_61_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[42]_reg  (.CLK(clknet_leaf_57_clk_i_regs),
    .RESET_B(net1529),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_036_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_364_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2026]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[43]_reg  (.CLK(clknet_leaf_61_clk_i_regs),
    .RESET_B(net1528),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_037_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_363_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2027]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[44]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_038_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2028]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_362_ ),
    .CLK(clknet_leaf_51_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[45]_reg  (.RESET_B(net1589),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_039_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2029]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_361_ ),
    .CLK(clknet_leaf_52_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[46]_reg  (.CLK(clknet_leaf_52_clk_i_regs),
    .RESET_B(net1589),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_040_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_360_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2030]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[47]_reg  (.CLK(clknet_leaf_52_clk_i_regs),
    .RESET_B(net1589),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_041_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_359_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2031]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[48]_reg  (.RESET_B(net1587),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_042_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2032]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_358_ ),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[49]_reg  (.CLK(clknet_leaf_13_clk_i_regs),
    .RESET_B(net1587),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_043_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_357_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2033]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[4]_reg  (.CLK(clknet_leaf_65_clk_i_regs),
    .RESET_B(net1534),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_044_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_356_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1988]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[50]_reg  (.RESET_B(net1616),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_045_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2034]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_355_ ),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[51]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1616),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_046_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_354_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2035]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[52]_reg  (.RESET_B(net1616),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_047_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2036]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_353_ ),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[53]_reg  (.RESET_B(net1616),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_048_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2037]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_352_ ),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[54]_reg  (.RESET_B(net1614),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_049_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2038]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_351_ ),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[55]_reg  (.CLK(clknet_leaf_11_clk_i_regs),
    .RESET_B(net1615),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_050_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_350_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2039]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[56]_reg  (.CLK(clknet_leaf_13_clk_i_regs),
    .RESET_B(net1615),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_051_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_349_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2040]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[57]_reg  (.CLK(clknet_leaf_12_clk_i_regs),
    .RESET_B(net1584),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_052_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_348_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2041]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[58]_reg  (.CLK(clknet_leaf_11_clk_i_regs),
    .RESET_B(net1614),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_053_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_347_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2042]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[59]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_054_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2043]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_346_ ),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[5]_reg  (.CLK(clknet_leaf_59_clk_i_regs),
    .RESET_B(net1528),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_055_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_345_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1989]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[60]_reg  (.CLK(clknet_leaf_11_clk_i_regs),
    .RESET_B(net1584),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_056_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_344_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2044]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[61]_reg  (.CLK(clknet_leaf_12_clk_i_regs),
    .RESET_B(net1585),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_057_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_343_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2045]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[62]_reg  (.CLK(clknet_leaf_12_clk_i_regs),
    .RESET_B(net1615),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_058_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_342_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2046]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[63]_reg  (.CLK(clknet_leaf_12_clk_i_regs),
    .RESET_B(net1585),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_059_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_341_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [2047]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[6]_reg  (.RESET_B(net1529),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_060_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1990]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_340_ ),
    .CLK(clknet_leaf_59_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[7]_reg  (.RESET_B(net1529),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_061_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1991]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_339_ ),
    .CLK(clknet_leaf_57_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[8]_reg  (.RESET_B(net1530),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_062_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1992]),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_338_ ),
    .CLK(clknet_leaf_55_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/mcycle_counter_i/counter_val_o[9]_reg  (.CLK(clknet_leaf_57_clk_i_regs),
    .RESET_B(net1528),
    .D(\i_ibex/cs_registers_i/mcycle_counter_i/_063_ ),
    .Q_N(\i_ibex/cs_registers_i/mcycle_counter_i/_337_ ),
    .Q(\i_ibex/cs_registers_i/mhpmcounter [1993]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0522_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0064_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [62]),
    .VSS(VSS));
 sg13g2_buf_2 fanout908 (.A(net909),
    .X(net908),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0524_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [24]),
    .B(\i_ibex/cs_registers_i/minstret_raw [25]),
    .C(\i_ibex/cs_registers_i/minstret_raw [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(net910),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0526_  (.A(\i_ibex/cs_registers_i/minstret_raw [27]),
    .B(\i_ibex/cs_registers_i/minstret_raw [28]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0527_  (.A(\i_ibex/cs_registers_i/minstret_raw [29]),
    .B(\i_ibex/cs_registers_i/minstret_raw [30]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0068_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0528_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0070_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [31]),
    .VSS(VSS));
 sg13g2_buf_2 fanout906 (.A(\i_ibex/cs_registers_i/dscratch1_en ),
    .X(net906),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0530_  (.B(net1492),
    .C(\i_ibex/cs_registers_i/minstret_raw [18]),
    .A(net1493),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0072_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_raw [19]));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0533_  (.B(\i_ibex/cs_registers_i/minstret_raw [21]),
    .C(\i_ibex/cs_registers_i/minstret_raw [22]),
    .A(\i_ibex/cs_registers_i/minstret_raw [20]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0075_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_raw [23]));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0534_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0070_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0072_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0075_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0535_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout903 (.X(net903),
    .A(net905),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0537_  (.A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .B(\i_ibex/cs_registers_i/minstret_raw [41]),
    .C(\i_ibex/cs_registers_i/minstret_raw [42]),
    .D(\i_ibex/cs_registers_i/minstret_raw [43]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0538_  (.A(\i_ibex/cs_registers_i/minstret_raw [44]),
    .B(\i_ibex/cs_registers_i/minstret_raw [45]),
    .C(\i_ibex/cs_registers_i/minstret_raw [46]),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0079_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(net905),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0540_  (.B(\i_ibex/cs_registers_i/minstret_raw [33]),
    .C(\i_ibex/cs_registers_i/minstret_raw [34]),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0541_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0083_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [38]),
    .B(\i_ibex/cs_registers_i/minstret_raw [39]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout901 (.X(net901),
    .A(net906),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0543_  (.B(\i_ibex/cs_registers_i/minstret_raw [36]),
    .C(\i_ibex/cs_registers_i/minstret_raw [37]),
    .A(\i_ibex/cs_registers_i/minstret_raw [35]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0085_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(\i_ibex/cs_registers_i/mie_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0545_  (.B(\i_ibex/cs_registers_i/minstret_raw [15]),
    .C(\i_ibex/cs_registers_i/minstret_raw [47]),
    .A(\i_ibex/cs_registers_i/minstret_raw [14]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0087_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0546_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0082_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0083_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0085_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0088_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0087_ ));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0547_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0089_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [7]),
    .B(\i_ibex/cs_registers_i/minstret_raw [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0548_  (.B(\i_ibex/cs_registers_i/minstret_raw [11]),
    .C(\i_ibex/cs_registers_i/minstret_raw [9]),
    .A(\i_ibex/cs_registers_i/minstret_raw [10]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0090_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout899 (.A(net900),
    .X(net899),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0550_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0092_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [0]),
    .B(\i_ibex/cs_registers_i/minstret_raw [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0551_  (.B(\i_ibex/cs_registers_i/minstret_raw [3]),
    .C(\i_ibex/cs_registers_i/minstret_raw [4]),
    .A(\i_ibex/cs_registers_i/minstret_raw [2]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0552_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0089_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0090_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0092_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0094_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0093_ ));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(net900),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0554_  (.A(\i_ibex/cs_registers_i/minstret_raw [12]),
    .B(\i_ibex/cs_registers_i/minstret_raw [13]),
    .C(\i_ibex/cs_registers_i/minstret_raw [5]),
    .D(\i_ibex/cs_registers_i/minstret_raw [6]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0096_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0555_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0088_ ),
    .C(net693),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0080_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0096_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0556_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0098_ ),
    .B(net1397),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(\i_ibex/cs_registers_i/mtvec_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0558_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0100_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [56]),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0559_  (.B(\i_ibex/cs_registers_i/minstret_raw [52]),
    .C(\i_ibex/cs_registers_i/minstret_raw [53]),
    .A(\i_ibex/cs_registers_i/minstret_raw [51]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0560_  (.B(\i_ibex/cs_registers_i/minstret_raw [49]),
    .C(\i_ibex/cs_registers_i/minstret_raw [50]),
    .A(\i_ibex/cs_registers_i/minstret_raw [48]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(\i_ibex/cs_registers_i/mtvec_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0562_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0104_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [54]),
    .B(\i_ibex/cs_registers_i/minstret_raw [55]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0563_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0100_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0101_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0102_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0104_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0564_  (.A(\i_ibex/cs_registers_i/minstret_raw [57]),
    .B(\i_ibex/cs_registers_i/minstret_raw [58]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0565_  (.A(\i_ibex/cs_registers_i/minstret_raw [60]),
    .B(\i_ibex/cs_registers_i/minstret_raw [61]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0107_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0566_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0105_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0106_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [59]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0108_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0107_ ));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0567_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0064_ ),
    .B(net1386),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0108_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0109_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0568_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0109_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [63]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [63]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(net896),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0570_  (.A(net1387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0108_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0571_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [62]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0064_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0572_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0112_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [52]),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0573_  (.B(\i_ibex/cs_registers_i/minstret_raw [49]),
    .C(\i_ibex/cs_registers_i/minstret_raw [50]),
    .A(\i_ibex/cs_registers_i/minstret_raw [48]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0113_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_raw [51]));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0574_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0114_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0113_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0112_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0575_  (.A(net1386),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0114_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0576_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0115_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [53]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [53]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0577_  (.A(net1386),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0113_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0578_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [52]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0112_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0579_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0098_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0102_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0117_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0580_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0117_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [51]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [51]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0581_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0118_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [48]),
    .B(\i_ibex/cs_registers_i/minstret_raw [49]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0582_  (.A(net1386),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0118_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0583_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0119_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [50]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [50]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0584_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0120_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [48]),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0585_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0120_ ),
    .B(net1386),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0586_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0121_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [49]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [49]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0587_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [48]),
    .A(\i_ibex/cs_registers_i/minstret_raw [48]),
    .B(net1386),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0588_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0082_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0083_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0085_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/cs_registers_i/minstret_counter_i/_0589_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0590_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [14]),
    .B(\i_ibex/cs_registers_i/minstret_raw [15]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0096_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(\i_ibex/cs_registers_i/mtvec_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0592_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0076_ ),
    .C(net693),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0126_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net894),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0594_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0126_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0595_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0129_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0080_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0596_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [47]),
    .A(\i_ibex/cs_registers_i/minstret_raw [47]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0597_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0130_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [44]),
    .B(\i_ibex/cs_registers_i/minstret_raw [45]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0598_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0131_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0130_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0599_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [46]),
    .A(\i_ibex/cs_registers_i/minstret_raw [46]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0600_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0132_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [44]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0601_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .B(net1385),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0132_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0602_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0133_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [45]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [45]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0603_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0134_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0079_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0604_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [44]),
    .A(\i_ibex/cs_registers_i/minstret_raw [44]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0134_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0605_  (.B(\i_ibex/cs_registers_i/minstret_raw [60]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0105_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [59]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0135_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0106_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0606_  (.A(net1387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0135_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0607_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0136_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [61]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [61]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0608_  (.B(\i_ibex/cs_registers_i/minstret_raw [41]),
    .C(\i_ibex/cs_registers_i/minstret_raw [42]),
    .A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0609_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0137_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .C(net1385),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0138_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0610_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0138_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [43]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [43]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0611_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0139_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .B(\i_ibex/cs_registers_i/minstret_raw [41]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0612_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0139_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .C(net1385),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0140_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0613_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0140_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [42]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [42]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0614_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0141_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0615_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [41]),
    .A(\i_ibex/cs_registers_i/minstret_raw [41]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0616_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0128_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [40]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0617_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0142_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0082_ ),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0618_  (.B(\i_ibex/cs_registers_i/minstret_raw [36]),
    .C(\i_ibex/cs_registers_i/minstret_raw [37]),
    .A(\i_ibex/cs_registers_i/minstret_raw [35]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0143_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0142_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0619_  (.A(net1385),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0143_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0620_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0145_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [38]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0621_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [39]),
    .A(\i_ibex/cs_registers_i/minstret_raw [39]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0622_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0146_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [38]),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0623_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [38]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0146_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0624_  (.B(\i_ibex/cs_registers_i/minstret_raw [36]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0142_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [35]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0625_  (.A(net1385),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0147_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0148_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0626_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0148_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [37]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [37]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0627_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0149_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [35]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0628_  (.A(net1385),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0149_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0629_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0150_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [36]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [36]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0630_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0082_ ),
    .B(net1385),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0151_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0631_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0151_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [35]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [35]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0632_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0152_ ),
    .A(net693),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0633_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ),
    .B(net1384),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0153_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0634_  (.B(\i_ibex/cs_registers_i/minstret_raw [33]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0153_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0635_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [34]),
    .A(\i_ibex/cs_registers_i/minstret_raw [34]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0636_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0105_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0106_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [59]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0637_  (.A(net1386),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0155_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0156_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0638_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0156_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [60]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [60]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0639_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0157_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0153_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0640_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [33]),
    .A(\i_ibex/cs_registers_i/minstret_raw [33]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0641_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [32]),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .B(net1385),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0642_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0072_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0075_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0643_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0158_ ),
    .B(net693),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout892 (.A(\i_ibex/cs_registers_i/dscratch0_en ),
    .X(net892),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0645_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0161_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0646_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [31]),
    .A(\i_ibex/cs_registers_i/minstret_raw [31]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0647_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0162_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [29]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0648_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0163_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0162_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0649_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [30]),
    .A(\i_ibex/cs_registers_i/minstret_raw [30]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0650_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0164_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [28]),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0651_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [27]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0652_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0166_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0165_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0164_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0653_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [29]),
    .A(\i_ibex/cs_registers_i/minstret_raw [29]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0166_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0654_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [28]),
    .A(\i_ibex/cs_registers_i/minstret_raw [28]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0655_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0167_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0656_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [27]),
    .A(\i_ibex/cs_registers_i/minstret_raw [27]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0657_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0168_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [24]),
    .B(\i_ibex/cs_registers_i/minstret_raw [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/minstret_counter_i/_0658_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0169_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .A_N(\i_ibex/cs_registers_i/minstret_counter_i/_0168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0659_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [26]),
    .A(\i_ibex/cs_registers_i/minstret_raw [26]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0660_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0170_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [24]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0661_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [25]),
    .A(\i_ibex/cs_registers_i/minstret_raw [25]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0170_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0662_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [24]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0663_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0171_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0105_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0664_  (.A(net1386),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0171_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0172_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0665_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0172_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [59]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [59]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0666_  (.B(\i_ibex/cs_registers_i/minstret_raw [21]),
    .C(\i_ibex/cs_registers_i/minstret_raw [22]),
    .A(net1491),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0173_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout891 (.X(net891),
    .A(net892),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0668_  (.A(net1494),
    .B(net1492),
    .C(\i_ibex/cs_registers_i/minstret_raw [18]),
    .D(\i_ibex/cs_registers_i/minstret_raw [19]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0669_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0175_ ),
    .B(net693),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/minstret_counter_i/_0670_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0177_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .A_N(\i_ibex/cs_registers_i/minstret_counter_i/_0173_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0671_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [23]),
    .A(\i_ibex/cs_registers_i/minstret_raw [23]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0177_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0672_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0178_ ),
    .A(net1491),
    .B(\i_ibex/cs_registers_i/minstret_raw [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/minstret_counter_i/_0673_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0179_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .A_N(\i_ibex/cs_registers_i/minstret_counter_i/_0178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0674_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [22]),
    .A(\i_ibex/cs_registers_i/minstret_raw [22]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0179_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0675_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0180_ ),
    .A(net1491),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0676_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [21]),
    .A(\i_ibex/cs_registers_i/minstret_raw [21]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0180_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0677_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .A(net1491),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0678_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0181_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [18]),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0679_  (.A(net693),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0182_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0680_  (.B(net1492),
    .C(net1382),
    .A(net1494),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0183_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0681_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0184_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0183_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0181_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0682_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [19]),
    .A(\i_ibex/cs_registers_i/minstret_raw [19]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0683_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [18]),
    .A(\i_ibex/cs_registers_i/minstret_raw [18]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0183_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout890 (.A(\i_ibex/cs_registers_i/gen_trigger_regs.tmatch_value_we ),
    .X(net890),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0685_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0186_ ),
    .A(net1493),
    .B(net1383),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0686_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [17]),
    .A(net1492),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0186_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0687_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [16]),
    .A(net1494),
    .B(net1384),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0688_  (.A(net693),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0096_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0689_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0188_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [14]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0690_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [15]),
    .A(\i_ibex/cs_registers_i/minstret_raw [15]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0691_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0189_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [14]),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0692_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [14]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0189_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0693_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0190_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [57]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0694_  (.A(net1387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0190_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0191_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0695_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0191_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [58]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [58]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0696_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0089_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0090_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0697_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0193_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [5]),
    .B(\i_ibex/cs_registers_i/minstret_raw [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0698_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0092_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0093_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0193_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0699_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0192_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [12]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0195_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0700_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [13]),
    .A(\i_ibex/cs_registers_i/minstret_raw [13]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0195_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0701_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0089_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0092_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0093_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0196_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0193_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0702_  (.A(\i_ibex/cs_registers_i/minstret_raw [9]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0196_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0703_  (.B(\i_ibex/cs_registers_i/minstret_raw [11]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0197_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [10]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0704_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [12]),
    .A(\i_ibex/cs_registers_i/minstret_raw [12]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0705_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0199_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [10]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0706_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [11]),
    .A(\i_ibex/cs_registers_i/minstret_raw [11]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0199_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0707_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0200_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [10]),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0708_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [10]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0200_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0709_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0201_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [9]),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0710_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [9]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0201_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0711_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0092_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0093_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0712_  (.B(\i_ibex/cs_registers_i/minstret_raw [6]),
    .C(\i_ibex/cs_registers_i/minstret_raw [7]),
    .A(\i_ibex/cs_registers_i/minstret_raw [5]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0203_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0202_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0713_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [8]),
    .A(\i_ibex/cs_registers_i/minstret_raw [8]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0714_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [7]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0715_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0204_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [5]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0716_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [6]),
    .A(\i_ibex/cs_registers_i/minstret_raw [6]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0717_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0205_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [5]),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0718_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [5]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0205_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0719_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0206_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [3]),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0720_  (.B(\i_ibex/cs_registers_i/minstret_raw [1]),
    .C(\i_ibex/cs_registers_i/minstret_raw [2]),
    .A(\i_ibex/cs_registers_i/minstret_raw [0]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0721_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0208_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0207_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0206_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0722_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [4]),
    .A(\i_ibex/cs_registers_i/minstret_raw [4]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0208_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0723_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0101_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0102_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0724_  (.B(\i_ibex/cs_registers_i/minstret_raw [55]),
    .C(\i_ibex/cs_registers_i/minstret_raw [56]),
    .A(\i_ibex/cs_registers_i/minstret_raw [54]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0210_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0209_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0725_  (.A(net1387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0210_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0726_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0211_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [57]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [57]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0727_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [3]),
    .A(\i_ibex/cs_registers_i/minstret_raw [3]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0728_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [2]),
    .A(\i_ibex/cs_registers_i/minstret_raw [2]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0729_  (.B(\i_ibex/cs_registers_i/minstret_raw [1]),
    .A(\i_ibex/cs_registers_i/minstret_raw [0]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0730_  (.B(\i_ibex/cs_registers_i/minstret_raw [55]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0209_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [54]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0212_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0731_  (.A(net1387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0212_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0213_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0732_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [56]),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0100_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0213_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0733_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0214_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [54]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0734_  (.A(net1387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0214_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0215_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0735_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0215_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [55]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [55]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/cs_registers_i/minstret_counter_i/_0736_  (.A(net1387),
    .B_N(\i_ibex/cs_registers_i/minstret_counter_i/_0209_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0737_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0216_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [54]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [54]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(net890),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout888 (.A(net890),
    .X(net888),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout887 (.X(net887),
    .A(net888),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout886 (.A(net890),
    .X(net886),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(net890),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/cs_registers_i/minstret_counter_i/_0743_  (.A(net878),
    .B_N(net408),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0222_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0744_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0223_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0222_ ),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [0]),
    .A2(net878),
    .A1(net973),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(\i_ibex/cs_registers_i/mepc_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(net884),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_8 \i_ibex/cs_registers_i/minstret_counter_i/_0747_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0226_ ),
    .A(net390),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout882 (.A(net883),
    .X(net882),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0749_  (.B1(net387),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0228_ ),
    .VSS(VSS),
    .A1(net408),
    .A2(net878));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0750_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0229_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [0]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0751_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0229_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0000_ ),
    .VSS(VSS),
    .A1(net392),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0223_ ));
 sg13g2_buf_4 fanout881 (.X(net881),
    .A(\i_ibex/cs_registers_i/mepc_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout880 (.X(net880),
    .A(net881),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0754_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0232_ ),
    .A(net388),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0755_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0233_ ),
    .A(net410),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0756_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0232_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0200_ ),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0233_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout879 (.A(\i_ibex/cs_registers_i/mhpmcounter_we [2]),
    .X(net879),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0758_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0236_ ),
    .A(net877),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0759_  (.A(net390),
    .B(net846),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout878 (.X(net878),
    .A(net879),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout877 (.A(net879),
    .X(net877),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0762_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0240_ ),
    .B1(net828),
    .B2(net935),
    .A2(\i_ibex/cs_registers_i/minstret_raw [10]),
    .A1(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0763_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0240_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0001_ ),
    .VSS(VSS),
    .A1(net877),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0234_ ));
 sg13g2_and4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0764_  (.A(net408),
    .B(\i_ibex/cs_registers_i/minstret_raw [10]),
    .C(\i_ibex/cs_registers_i/minstret_raw [9]),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0196_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0241_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0765_  (.A(\i_ibex/cs_registers_i/minstret_raw [11]),
    .B(net876),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0766_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0243_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0241_ ),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0242_ ),
    .A2(net876),
    .A1(net937),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0767_  (.B1(net388),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0244_ ),
    .VSS(VSS),
    .A1(net876),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0241_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0768_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0245_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [11]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0769_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0245_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0002_ ),
    .VSS(VSS),
    .A1(net392),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0243_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0770_  (.A(net390),
    .B(\i_ibex/cs_registers_i/minstret_raw [12]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0771_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0192_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ),
    .A(net409),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0772_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0246_ ),
    .A1(\i_ibex/cs_registers_i/minstret_raw [12]),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0247_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0248_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0773_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0249_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0248_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0774_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0250_ ),
    .B1(net828),
    .B2(net939),
    .A2(\i_ibex/cs_registers_i/minstret_raw [12]),
    .A1(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0775_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0250_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0003_ ),
    .VSS(VSS),
    .A1(net876),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0249_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0776_  (.A(net390),
    .B(\i_ibex/cs_registers_i/minstret_raw [13]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0777_  (.B(\i_ibex/cs_registers_i/minstret_raw [12]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0192_ ),
    .A(net409),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0252_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0778_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0251_ ),
    .A1(\i_ibex/cs_registers_i/minstret_raw [13]),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0252_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0779_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0254_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0253_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0780_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0255_ ),
    .B1(net828),
    .B2(net957),
    .A2(\i_ibex/cs_registers_i/minstret_raw [13]),
    .A1(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0781_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0255_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0004_ ),
    .VSS(VSS),
    .A1(net879),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0254_ ));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0783_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net410),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0257_ ),
    .B1(\i_ibex/cs_registers_i/minstret_raw [14]));
 sg13g2_and4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0784_  (.A(net408),
    .B(net387),
    .C(\i_ibex/cs_registers_i/minstret_raw [14]),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0785_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0259_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0258_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0257_ ));
 sg13g2_nand2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0786_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0260_ ),
    .A(net387),
    .B(net877),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout875 (.A(\i_ibex/cs_registers_i/mscratch_en ),
    .X(net875),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0788_  (.A(net940),
    .B(net824),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0789_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0259_ ),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0262_ ),
    .B1(net846),
    .A1(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0005_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0189_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0790_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0263_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [14]),
    .B(\i_ibex/cs_registers_i/minstret_raw [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0791_  (.A(net383),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0222_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0792_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0264_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0265_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0793_  (.A(\i_ibex/cs_registers_i/minstret_raw [15]),
    .B(net824),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0794_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0187_ ),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0266_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0264_ ),
    .A1(net959),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0267_ ),
    .A2(net828));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0795_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0263_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0265_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0006_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0267_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0796_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0268_ ),
    .A(net410),
    .B(net1382),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0797_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0269_ ),
    .A(net408),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0798_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0269_ ),
    .B(net391),
    .C(net1493),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0152_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0270_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0799_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1493),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0268_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0271_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0270_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0800_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0272_ ),
    .B1(net828),
    .B2(net942),
    .A2(net1493),
    .A1(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0801_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0272_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0007_ ),
    .VSS(VSS),
    .A1(net878),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0271_ ));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0802_  (.B(net1492),
    .A(net1493),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0273_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0803_  (.A0(net943),
    .A1(net1492),
    .S(net824),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0804_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0275_ ),
    .A(net1382),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0805_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0273_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0274_ ),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0275_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0806_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0276_ ),
    .A(net387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0181_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0807_  (.B(net1493),
    .C(net1492),
    .A(net410),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0277_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net1382));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0808_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0276_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0181_ ),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0277_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0809_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0279_ ),
    .B1(net827),
    .B2(net946),
    .A2(\i_ibex/cs_registers_i/minstret_raw [18]),
    .A1(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0810_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0279_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0009_ ),
    .VSS(VSS),
    .A1(net879),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0278_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0811_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0280_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [19]),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0812_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0281_ ),
    .A(net408),
    .B(net1492),
    .C(\i_ibex/cs_registers_i/minstret_raw [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0813_  (.B(net693),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .A(net1493),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0282_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0281_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0814_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net847),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0282_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0283_ ),
    .B1(net392));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0816_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0285_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0280_ ),
    .B(net847),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0817_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0286_ ),
    .A(net948),
    .B(net878),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0818_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0286_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0287_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0282_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0285_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0819_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0288_ ),
    .A(net389),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0287_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0820_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0288_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0010_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0280_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0283_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0821_  (.B(\i_ibex/cs_registers_i/minstret_raw [0]),
    .C(\i_ibex/cs_registers_i/minstret_raw [1]),
    .A(net408),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0289_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0822_  (.A0(net971),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0289_ ),
    .S(net846),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0290_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0823_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net410),
    .A2(\i_ibex/cs_registers_i/minstret_raw [0]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0291_ ),
    .B1(net876));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0824_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0292_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [1]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0825_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0292_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0293_ ),
    .VSS(VSS),
    .A1(net391),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0291_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0826_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0293_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0294_ ),
    .VSS(VSS),
    .A1(net392),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0290_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0827_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0011_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0294_ ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0828_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0295_ ),
    .A(net409),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0829_  (.A(net390),
    .B(net1491),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0830_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0297_ ),
    .A(net408),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0176_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0831_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1491),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0295_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0298_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0297_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0832_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0299_ ),
    .B1(net827),
    .B2(net426),
    .A2(net1491),
    .A1(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0833_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0299_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0012_ ),
    .VSS(VSS),
    .A1(net879),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0298_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0834_  (.A(net961),
    .B(net827),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0835_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [21]),
    .A2(net825),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0301_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0300_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0836_  (.B(net1382),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0264_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0175_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0837_  (.B(\i_ibex/cs_registers_i/minstret_raw [21]),
    .A(net1491),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0838_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0303_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0304_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0839_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0301_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0013_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0304_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0840_  (.A(net412),
    .B(net826),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0841_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [22]),
    .A2(net825),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0306_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0305_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0842_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0307_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [22]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0843_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0307_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0308_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0844_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0306_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0014_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0308_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0845_  (.A(net414),
    .B(net826),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0309_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0846_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [23]),
    .A2(net825),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0310_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0309_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0847_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0311_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [23]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0173_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0848_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0311_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0849_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0302_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0310_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0015_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0312_ ));
 sg13g2_nor2_2 \i_ibex/cs_registers_i/minstret_counter_i/_0850_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0093_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0289_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0851_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0192_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0158_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0314_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0313_ ));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0852_  (.A(\i_ibex/cs_registers_i/minstret_raw [24]),
    .B(net878),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0314_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0853_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net928),
    .A2(net878),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0316_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0315_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0854_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net847),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0314_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0317_ ),
    .B1(net391));
 sg13g2_nand2b_1 \i_ibex/cs_registers_i/minstret_counter_i/_0855_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0318_ ),
    .B(\i_ibex/cs_registers_i/minstret_raw [24]),
    .A_N(\i_ibex/cs_registers_i/minstret_counter_i/_0317_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0856_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0318_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0016_ ),
    .VSS(VSS),
    .A1(net391),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0316_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0857_  (.A(net416),
    .B(net826),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0858_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [25]),
    .A2(net825),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0320_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0319_ ));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0859_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0094_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0124_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0158_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0264_ ));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0860_  (.B(\i_ibex/cs_registers_i/minstret_raw [25]),
    .A(\i_ibex/cs_registers_i/minstret_raw [24]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0861_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0322_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0862_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0320_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0017_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0323_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0863_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0324_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [26]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0864_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0325_ ),
    .A(net387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0324_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0865_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0168_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0314_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0326_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0866_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0324_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0325_ ),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0326_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0327_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0867_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0328_ ),
    .B1(net826),
    .B2(net930),
    .A2(\i_ibex/cs_registers_i/minstret_raw [26]),
    .A1(net392),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0868_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0328_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0018_ ),
    .VSS(VSS),
    .A1(net879),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0327_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0869_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0167_ ),
    .C(net825),
    .A(\i_ibex/cs_registers_i/minstret_raw [27]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0870_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0324_ ),
    .B(\i_ibex/cs_registers_i/minstret_raw [27]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0168_ ),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0871_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net424),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0330_ ),
    .B1(net826),
    .A1(\i_ibex/cs_registers_i/minstret_raw [27]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0331_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0228_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0872_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0019_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0329_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0331_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0873_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0332_ ),
    .A(net387),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0164_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0874_  (.B(\i_ibex/cs_registers_i/minstret_raw [27]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .A(net409),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0333_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0159_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0875_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0332_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0164_ ),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0333_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0334_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0876_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0335_ ),
    .B1(net826),
    .B2(net419),
    .A2(\i_ibex/cs_registers_i/minstret_raw [28]),
    .A1(net392),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0877_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0335_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0020_ ),
    .VSS(VSS),
    .A1(net878),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0334_ ));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0878_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0336_ ),
    .A(net420),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0879_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0337_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0880_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0338_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0066_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0881_  (.B1(net847),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0339_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0338_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0314_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0882_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net388),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0339_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0340_ ),
    .B1(\i_ibex/cs_registers_i/minstret_raw [29]));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0883_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0162_ ),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0340_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0337_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0336_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0021_ ),
    .A2(net826));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0884_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0341_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [2]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0885_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0342_ ),
    .A(net387),
    .B(\i_ibex/cs_registers_i/minstret_raw [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0886_  (.B(\i_ibex/cs_registers_i/minstret_raw [0]),
    .C(\i_ibex/cs_registers_i/minstret_raw [1]),
    .A(net409),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0887_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0344_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0341_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0888_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0344_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0345_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0342_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0343_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0889_  (.A(net949),
    .B(net824),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0346_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0890_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0345_ ),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0346_ ),
    .B1(net846),
    .A1(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0022_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0341_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0891_  (.A(net963),
    .B(net826),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0347_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0892_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [30]),
    .A2(net824),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0348_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0347_ ));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0893_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0162_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [30]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0349_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0894_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0349_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0350_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0895_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0348_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0023_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0350_ ));
 sg13g2_and2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0896_  (.A(net422),
    .B(net827),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0351_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0897_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [31]),
    .A2(net824),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0352_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0351_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0898_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0353_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0070_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0899_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0353_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0354_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0900_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0321_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0352_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0024_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0354_ ));
 sg13g2_and3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0901_  (.X(\i_ibex/cs_registers_i/minstret_counter_i/_0355_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0076_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0222_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout873 (.A(net874),
    .X(net873),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0903_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0357_ ),
    .A(net1383),
    .B(net823),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0904_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0358_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0357_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0905_  (.A0(net973),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0358_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0906_  (.B(net1383),
    .C(net823),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0359_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0907_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0360_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [33]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0359_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0908_  (.A0(net971),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0360_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0909_  (.B(\i_ibex/cs_registers_i/minstret_raw [33]),
    .C(net1383),
    .A(\i_ibex/cs_registers_i/minstret_raw [32]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0361_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net823));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0910_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0362_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [34]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0361_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0911_  (.A0(net949),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0362_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0912_  (.B(net1383),
    .C(net823),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0142_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0363_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0913_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0364_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [35]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0363_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(net873),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0915_  (.A0(net952),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0364_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0916_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0076_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0222_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0069_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0366_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(net875),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0918_  (.A(net1384),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0149_ ),
    .C(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0368_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0919_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0368_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [36]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0369_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0920_  (.A0(net953),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0369_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0921_  (.A(net1384),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0147_ ),
    .C(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0370_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0922_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0370_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [37]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0371_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0923_  (.A0(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0371_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0924_  (.A(net1384),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0143_ ),
    .C(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0925_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0373_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0146_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0926_  (.A0(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0373_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(net871),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0928_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0146_ ),
    .B(net1384),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0143_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0375_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net822));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0929_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0375_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [39]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0376_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0930_  (.A0(net955),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0376_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0931_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0377_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0207_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0269_ ));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0932_  (.A(net391),
    .B(\i_ibex/cs_registers_i/minstret_raw [3]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0377_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0378_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0933_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [3]),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0377_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0379_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0378_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0934_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0380_ ),
    .B1(net828),
    .B2(net952),
    .A2(\i_ibex/cs_registers_i/minstret_raw [3]),
    .A1(net392),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0935_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0380_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0033_ ),
    .VSS(VSS),
    .A1(net876),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0379_ ));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0936_  (.B(net1383),
    .C(net823),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0381_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0937_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0382_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0381_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0938_  (.A0(net931),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0382_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0939_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .C(net1383),
    .A(\i_ibex/cs_registers_i/minstret_raw [40]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0383_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net823));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0940_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0384_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [41]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0383_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0941_  (.A0(net933),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0384_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0942_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0139_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .C(net1384),
    .D(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0385_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0943_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0386_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [42]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0385_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0944_  (.A(net388),
    .B(net935),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0387_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0945_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net388),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0386_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0036_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0387_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0946_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0137_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .C(net1384),
    .D(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0388_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0947_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0388_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [43]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0389_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0948_  (.A0(net937),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0389_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0949_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .C(net1382),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0079_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0390_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0355_ ));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0950_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0391_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [44]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0951_  (.A0(net939),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0391_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0952_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0123_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0152_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0132_ ),
    .D(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0392_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0953_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0393_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [45]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0392_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0954_  (.A(net388),
    .B(net957),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0394_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0955_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net388),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0393_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0039_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0394_ ));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0956_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .C(net1382),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0130_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0395_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net823));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0957_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0396_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [46]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0395_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0958_  (.A0(net940),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0396_ ),
    .S(net384),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0959_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0122_ ),
    .C(net1382),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0080_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0397_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net823));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0960_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0398_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [47]),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(\i_ibex/cs_registers_i/mtval_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0962_  (.A0(net959),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0398_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(net869),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0964_  (.A(net1397),
    .B(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0401_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0965_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0402_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0120_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0401_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0966_  (.A0(net941),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0402_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0967_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0120_ ),
    .B(net1397),
    .C(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0403_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0968_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0403_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [49]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0404_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0969_  (.A0(net943),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0404_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0970_  (.B1(\i_ibex/cs_registers_i/minstret_raw [4]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0405_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0206_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0377_ ));
 sg13g2_or4_1 \i_ibex/cs_registers_i/minstret_counter_i/_0971_  (.A(net393),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0206_ ),
    .C(\i_ibex/cs_registers_i/minstret_raw [4]),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0377_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0406_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0972_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0407_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0405_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0406_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_0973_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0408_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0407_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_0974_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0409_ ),
    .B1(net828),
    .B2(net953),
    .A2(\i_ibex/cs_registers_i/minstret_raw [4]),
    .A1(net392),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_0975_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0409_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0044_ ),
    .VSS(VSS),
    .A1(net876),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0408_ ));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0976_  (.A(net1397),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0118_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0410_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0977_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0410_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [50]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0411_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0978_  (.A0(net946),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0411_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0979_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0097_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0102_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0412_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0980_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0412_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [51]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0413_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0981_  (.A0(net948),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0413_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0982_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0097_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0113_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0414_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0983_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0415_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0112_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0414_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0984_  (.A0(net427),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0415_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0985_  (.A(net1397),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0114_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0416_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0986_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0416_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [53]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0417_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0987_  (.A0(net961),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0417_ ),
    .S(net386),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/cs_registers_i/minstret_counter_i/_0988_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0101_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0102_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0418_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net820));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0989_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0418_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [54]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0419_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0990_  (.A0(net412),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0419_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0991_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0214_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0420_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0992_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0420_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [55]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0421_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0993_  (.A0(net414),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0421_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_0994_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0212_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0422_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0995_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0423_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0100_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0422_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0996_  (.A0(net927),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0423_ ),
    .S(net385),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_0997_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0210_ ),
    .C(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0424_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0998_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0424_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [57]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0425_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_0999_  (.A0(net416),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0425_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1000_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0190_ ),
    .C(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0426_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1001_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0426_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [58]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0427_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1002_  (.A0(net930),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0427_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1003_  (.A(net1397),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0171_ ),
    .C(net822),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0428_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1004_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0428_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [59]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0429_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1005_  (.A0(net425),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0429_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1006_  (.B(net846),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0313_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [5]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0430_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_1007_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0430_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0431_ ),
    .VSS(VSS),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .A2(net846));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_1008_  (.B1(net388),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0432_ ),
    .VSS(VSS),
    .A1(net877),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0313_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1009_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0055_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0432_ ),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0205_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0431_ ),
    .A1(net387),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/cs_registers_i/minstret_counter_i/_1010_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0155_ ),
    .C(net820),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0433_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1011_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0433_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [60]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0434_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1012_  (.A0(net418),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0434_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1013_  (.A(net1397),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0135_ ),
    .C(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0435_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1014_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0435_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [61]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0436_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1015_  (.A0(net421),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0436_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1016_  (.A(net1398),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0108_ ),
    .C(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0437_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1017_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0438_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0064_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0437_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1018_  (.A0(net963),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0438_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0058_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_1019_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0064_ ),
    .B(net1397),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0108_ ),
    .D(net821),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0439_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1020_  (.B(\i_ibex/cs_registers_i/minstret_counter_i/_0439_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [63]),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0440_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1021_  (.A0(net422),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0440_ ),
    .S(net383),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/cs_registers_i/minstret_counter_i/_1022_  (.VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0441_ ),
    .A(\i_ibex/cs_registers_i/minstret_raw [6]),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1023_  (.B(\i_ibex/cs_registers_i/minstret_raw [5]),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0202_ ),
    .A(net409),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0442_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1024_  (.A(net390),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0441_ ),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0442_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0443_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/cs_registers_i/minstret_counter_i/_1025_  (.A2(\i_ibex/cs_registers_i/minstret_counter_i/_0442_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0441_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0443_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0444_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1026_  (.A(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .B(net824),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0445_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1027_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0444_ ),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0445_ ),
    .B1(net846),
    .A1(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0060_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0441_ ));
 sg13g2_nand2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1028_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0446_ ),
    .A(net409),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/cs_registers_i/minstret_counter_i/_1029_  (.A(\i_ibex/cs_registers_i/minstret_raw [7]),
    .B(net877),
    .C(\i_ibex/cs_registers_i/minstret_counter_i/_0446_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0447_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1030_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net955),
    .A2(net877),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0448_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0447_ ));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1031_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net409),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0194_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0449_ ),
    .B1(net877));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_1032_  (.B1(\i_ibex/cs_registers_i/minstret_raw [7]),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0450_ ),
    .VSS(VSS),
    .A1(net391),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0449_ ));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_1033_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0450_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0061_ ),
    .VSS(VSS),
    .A1(net391),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0448_ ));
 sg13g2_or2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1034_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0451_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0203_ ),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0269_ ));
 sg13g2_nor4_1 \i_ibex/cs_registers_i/minstret_counter_i/_1035_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0269_ ),
    .B(net391),
    .C(\i_ibex/cs_registers_i/minstret_raw [8]),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0203_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0452_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1036_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/minstret_raw [8]),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0451_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0453_ ),
    .B1(\i_ibex/cs_registers_i/minstret_counter_i/_0452_ ));
 sg13g2_a22oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1037_  (.Y(\i_ibex/cs_registers_i/minstret_counter_i/_0454_ ),
    .B1(net828),
    .B2(net931),
    .A2(\i_ibex/cs_registers_i/minstret_raw [8]),
    .A1(net390),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/cs_registers_i/minstret_counter_i/_1038_  (.B1(\i_ibex/cs_registers_i/minstret_counter_i/_0454_ ),
    .VDD(VDD),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0062_ ),
    .VSS(VSS),
    .A1(net876),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0453_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1039_  (.A(net390),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0201_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0455_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1040_  (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0089_ ),
    .B(\i_ibex/cs_registers_i/minstret_counter_i/_0446_ ),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0456_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1041_  (.A0(\i_ibex/cs_registers_i/minstret_counter_i/_0201_ ),
    .A1(\i_ibex/cs_registers_i/minstret_counter_i/_0455_ ),
    .S(\i_ibex/cs_registers_i/minstret_counter_i/_0456_ ),
    .X(\i_ibex/cs_registers_i/minstret_counter_i/_0457_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/minstret_counter_i/_1042_  (.A(net933),
    .B(net824),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0458_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/cs_registers_i/minstret_counter_i/_1043_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/cs_registers_i/minstret_counter_i/_0457_ ),
    .C1(\i_ibex/cs_registers_i/minstret_counter_i/_0458_ ),
    .B1(net846),
    .A1(net393),
    .Y(\i_ibex/cs_registers_i/minstret_counter_i/_0063_ ),
    .A2(\i_ibex/cs_registers_i/minstret_counter_i/_0201_ ));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[0]_reg  (.RESET_B(net1588),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0000_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [0]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/counter_val_upd_o [0]),
    .CLK(clknet_leaf_54_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[10]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0001_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [10]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0521_ ),
    .CLK(clknet_leaf_55_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[11]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0002_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [11]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0520_ ),
    .CLK(clknet_leaf_55_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[12]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0003_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [12]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0519_ ),
    .CLK(clknet_leaf_55_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[13]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0004_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [13]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0518_ ),
    .CLK(clknet_leaf_54_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[14]_reg  (.RESET_B(net1588),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0005_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [14]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0517_ ),
    .CLK(clknet_leaf_54_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[15]_reg  (.RESET_B(net1588),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0006_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [15]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0516_ ),
    .CLK(clknet_leaf_53_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[16]_reg  (.CLK(clknet_leaf_53_clk_i_regs),
    .RESET_B(net1588),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0007_ ),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0515_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[17]_reg  (.CLK(clknet_leaf_17_clk_i_regs),
    .RESET_B(net1588),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0008_ ),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0514_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[18]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0009_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [18]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0513_ ),
    .CLK(clknet_leaf_53_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[19]_reg  (.RESET_B(net1588),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0010_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [19]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0512_ ),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[1]_reg  (.RESET_B(net1602),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0011_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [1]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0511_ ),
    .CLK(clknet_leaf_59_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[20]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0012_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [20]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0510_ ),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[21]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0013_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [21]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0509_ ),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[22]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0014_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [22]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0508_ ),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[23]_reg  (.RESET_B(net1586),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0015_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [23]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0507_ ),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[24]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0016_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [24]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0506_ ),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[25]_reg  (.RESET_B(net1585),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0017_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [25]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0505_ ),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[26]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0018_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [26]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0504_ ),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[27]_reg  (.RESET_B(net1623),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0019_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [27]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0503_ ),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[28]_reg  (.RESET_B(net1586),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0020_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [28]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0502_ ),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[29]_reg  (.RESET_B(net1586),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0021_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [29]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0501_ ),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[2]_reg  (.RESET_B(net1602),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0022_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [2]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0500_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[30]_reg  (.RESET_B(net1585),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0023_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [30]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0499_ ),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[31]_reg  (.RESET_B(net1588),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0024_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [31]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0498_ ),
    .CLK(clknet_leaf_54_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[32]_reg  (.RESET_B(net1534),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0025_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [32]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0497_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[33]_reg  (.RESET_B(net1534),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0026_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [33]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0496_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[34]_reg  (.RESET_B(net1534),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0027_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [34]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0495_ ),
    .CLK(clknet_leaf_65_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[35]_reg  (.RESET_B(net1608),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0028_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [35]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0494_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[36]_reg  (.RESET_B(net1608),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0029_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [36]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0493_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[37]_reg  (.RESET_B(net1608),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0030_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [37]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0492_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[38]_reg  (.RESET_B(net1535),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0031_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [38]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0491_ ),
    .CLK(clknet_leaf_67_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[39]_reg  (.RESET_B(net1535),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0032_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [39]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0490_ ),
    .CLK(clknet_leaf_67_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[3]_reg  (.RESET_B(net1602),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0033_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [3]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0489_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[40]_reg  (.RESET_B(net1528),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0034_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [40]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0488_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[41]_reg  (.RESET_B(net1528),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0035_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [41]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0487_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[42]_reg  (.RESET_B(net1601),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0036_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [42]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0486_ ),
    .CLK(clknet_leaf_57_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[43]_reg  (.RESET_B(net1528),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0037_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [43]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0485_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[44]_reg  (.RESET_B(net1530),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0038_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [44]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0484_ ),
    .CLK(clknet_leaf_56_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[45]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0039_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [45]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0483_ ),
    .CLK(clknet_leaf_54_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[46]_reg  (.RESET_B(net1591),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0040_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [46]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0482_ ),
    .CLK(clknet_leaf_52_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[47]_reg  (.RESET_B(net1588),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0041_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [47]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0481_ ),
    .CLK(clknet_leaf_53_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[48]_reg  (.RESET_B(net1637),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0042_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [48]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0480_ ),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[49]_reg  (.RESET_B(net1616),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0043_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [49]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0479_ ),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[4]_reg  (.RESET_B(net1602),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0044_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [4]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0478_ ),
    .CLK(clknet_leaf_66_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[50]_reg  (.RESET_B(net1637),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0045_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [50]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0477_ ),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[51]_reg  (.RESET_B(net1637),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0046_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [51]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0476_ ),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[52]_reg  (.CLK(clknet_leaf_8_clk_i_regs),
    .RESET_B(net1618),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0047_ ),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0475_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [52]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[53]_reg  (.RESET_B(net1618),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0048_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [53]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0474_ ),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[54]_reg  (.RESET_B(net1637),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0049_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [54]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0473_ ),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[55]_reg  (.RESET_B(net1637),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0050_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [55]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0472_ ),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[56]_reg  (.CLK(clknet_leaf_9_clk_i_regs),
    .RESET_B(net1641),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0051_ ),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0471_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [56]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[57]_reg  (.RESET_B(net1614),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0052_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [57]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0470_ ),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[58]_reg  (.RESET_B(net1614),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0053_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [58]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0469_ ),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[59]_reg  (.RESET_B(net1614),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0054_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [59]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0468_ ),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[5]_reg  (.RESET_B(net1602),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0055_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [5]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0467_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[60]_reg  (.RESET_B(net1615),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0056_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [60]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0466_ ),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[61]_reg  (.RESET_B(net1614),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0057_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [61]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0465_ ),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[62]_reg  (.CLK(clknet_leaf_9_clk_i_regs),
    .RESET_B(net1614),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0058_ ),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0464_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [62]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[63]_reg  (.RESET_B(net1614),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0059_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [63]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0463_ ),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[6]_reg  (.RESET_B(net1602),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0060_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [6]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0462_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[7]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0061_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [7]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0461_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[8]_reg  (.RESET_B(net1598),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0062_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [8]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0460_ ),
    .CLK(clknet_leaf_58_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/minstret_counter_i/counter_val_o[9]_reg  (.RESET_B(net1601),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/minstret_counter_i/_0063_ ),
    .Q(\i_ibex/cs_registers_i/minstret_raw [9]),
    .Q_N(\i_ibex/cs_registers_i/minstret_counter_i/_0459_ ),
    .CLK(clknet_leaf_57_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/priv_mode_id_o[0]_reg  (.CLK(clknet_leaf_75_clk_i_regs),
    .RESET_B(net1573),
    .D(\i_ibex/cs_registers_i/_0004_ ),
    .Q_N(\i_ibex/priv_mode_id [0]),
    .Q(\i_ibex/cs_registers_i/_0000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/priv_mode_id_o[1]_reg  (.CLK(clknet_leaf_75_clk_i_regs),
    .RESET_B(net1573),
    .D(\i_ibex/cs_registers_i/_0005_ ),
    .Q_N(\i_ibex/priv_mode_id [1]),
    .Q(\i_ibex/cs_registers_i/_0001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(net868),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout866 (.A(net869),
    .X(net866),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_074_  (.A(\i_ibex/cs_registers_i/u_dcsr_csr/_000_ ),
    .B(net851),
    .Y(\i_ibex/cs_registers_i/u_dcsr_csr/_035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_dcsr_csr/_075_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/dcsr_d [0]),
    .A2(net851),
    .Y(\i_ibex/cs_registers_i/u_dcsr_csr/_003_ ),
    .B1(\i_ibex/cs_registers_i/u_dcsr_csr/_035_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_076_  (.A0(\i_ibex/cs_registers_i/dcsr_q [10]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [10]),
    .S(net853),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_077_  (.A0(\i_ibex/cs_registers_i/dcsr_q [11]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [11]),
    .S(net851),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_078_  (.A0(\i_ibex/debug_ebreaku ),
    .A1(\i_ibex/cs_registers_i/dcsr_d [12]),
    .S(net852),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_079_  (.A0(\i_ibex/cs_registers_i/dcsr_q [13]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [13]),
    .S(net856),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_081_  (.A0(\i_ibex/cs_registers_i/dcsr_q [14]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [14]),
    .S(net853),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_082_  (.A0(\i_ibex/debug_ebreakm ),
    .A1(\i_ibex/cs_registers_i/dcsr_d [15]),
    .S(net852),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_083_  (.A0(\i_ibex/cs_registers_i/dcsr_q [16]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [16]),
    .S(net854),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_084_  (.A0(\i_ibex/cs_registers_i/dcsr_q [17]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [17]),
    .S(net854),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_085_  (.A0(\i_ibex/cs_registers_i/dcsr_q [18]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [18]),
    .S(net854),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_086_  (.A0(\i_ibex/cs_registers_i/dcsr_q [19]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [19]),
    .S(net854),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_087_  (.A(\i_ibex/cs_registers_i/u_dcsr_csr/_001_ ),
    .B(net851),
    .Y(\i_ibex/cs_registers_i/u_dcsr_csr/_037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_dcsr_csr/_088_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/dcsr_d [1]),
    .A2(net851),
    .Y(\i_ibex/cs_registers_i/u_dcsr_csr/_014_ ),
    .B1(\i_ibex/cs_registers_i/u_dcsr_csr/_037_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_089_  (.A0(\i_ibex/cs_registers_i/dcsr_q [20]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [20]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_090_  (.A0(\i_ibex/cs_registers_i/dcsr_q [21]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [21]),
    .S(net854),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_091_  (.A0(\i_ibex/cs_registers_i/dcsr_q [22]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [22]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_092_  (.A0(\i_ibex/cs_registers_i/dcsr_q [23]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [23]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(net866),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_094_  (.A0(\i_ibex/cs_registers_i/dcsr_q [24]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [24]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_095_  (.A0(\i_ibex/cs_registers_i/dcsr_q [25]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [25]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_096_  (.A0(\i_ibex/cs_registers_i/dcsr_q [26]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [26]),
    .S(net854),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_097_  (.A0(\i_ibex/cs_registers_i/dcsr_q [27]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [27]),
    .S(net853),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_098_  (.A0(\i_ibex/cs_registers_i/dcsr_q [28]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [28]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_099_  (.A0(\i_ibex/cs_registers_i/dcsr_q [29]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [29]),
    .S(net852),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_100_  (.A0(\i_ibex/debug_single_step ),
    .A1(\i_ibex/cs_registers_i/dcsr_d [2]),
    .S(net853),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_101_  (.A(\i_ibex/cs_registers_i/u_dcsr_csr/_002_ ),
    .B(net854),
    .Y(\i_ibex/cs_registers_i/u_dcsr_csr/_039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_dcsr_csr/_102_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/dcsr_d [30]),
    .A2(net854),
    .Y(\i_ibex/cs_registers_i/u_dcsr_csr/_026_ ),
    .B1(\i_ibex/cs_registers_i/u_dcsr_csr/_039_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_103_  (.A0(\i_ibex/cs_registers_i/dcsr_q [31]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [31]),
    .S(net855),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_104_  (.A0(\i_ibex/cs_registers_i/dcsr_q [3]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [3]),
    .S(net851),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_105_  (.A0(\i_ibex/cs_registers_i/dcsr_q [4]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [4]),
    .S(net851),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_106_  (.A0(\i_ibex/cs_registers_i/dcsr_q [5]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [5]),
    .S(net851),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_107_  (.A0(\i_ibex/cs_registers_i/dcsr_q [6]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [6]),
    .S(net856),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_108_  (.A0(\i_ibex/cs_registers_i/dcsr_q [7]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [7]),
    .S(net852),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_109_  (.A0(\i_ibex/cs_registers_i/dcsr_q [8]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [8]),
    .S(net856),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dcsr_csr/_110_  (.A0(\i_ibex/cs_registers_i/dcsr_q [9]),
    .A1(\i_ibex/cs_registers_i/dcsr_d [9]),
    .S(net853),
    .X(\i_ibex/cs_registers_i/u_dcsr_csr/_034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1441__67  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net67));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1540),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/dcsr_q [0]),
    .Q(\i_ibex/cs_registers_i/u_dcsr_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1609),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_004_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_070_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_71_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_069_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_76_clk_i_regs),
    .RESET_B(net1542),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_068_ ),
    .Q(\i_ibex/debug_ebreaku ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1636),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_067_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1608),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[15]_reg  (.RESET_B(net1542),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_009_ ),
    .Q(\i_ibex/debug_ebreakm ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_065_ ),
    .CLK(clknet_leaf_76_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_064_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_4_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_063_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/dcsr_q [1]),
    .Q(\i_ibex/cs_registers_i/u_dcsr_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_1_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1640),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_8_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_1_clk_i_regs),
    .RESET_B(net1637),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_056_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_1_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1609),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_053_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_8_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_052_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_71_clk_i_regs),
    .RESET_B(net1608),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[2]_reg  (.RESET_B(net1609),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_025_ ),
    .Q(\i_ibex/debug_single_step ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_050_ ),
    .CLK(clknet_leaf_72_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[30]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/dcsr_q [30]),
    .Q(\i_ibex/cs_registers_i/u_dcsr_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_8_clk_i_regs),
    .RESET_B(net1616),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_049_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1542),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1542),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_047_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_71_clk_i_regs),
    .RESET_B(net1542),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_046_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[6]_reg  (.RESET_B(net1497),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_031_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [6]),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_045_ ),
    .CLK(clknet_leaf_76_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[7]_reg  (.RESET_B(net1542),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_032_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [7]),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_044_ ),
    .CLK(clknet_leaf_72_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[8]_reg  (.RESET_B(net1609),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_033_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [8]),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_043_ ),
    .CLK(clknet_leaf_72_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dcsr_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_70_clk_i_regs),
    .RESET_B(net1609),
    .D(\i_ibex/cs_registers_i/u_dcsr_csr/_034_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dcsr_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/dcsr_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout863 (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_087_ ),
    .X(net863),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_095_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_071_  (.A0(\i_ibex/csr_depc [0]),
    .A1(\i_ibex/cs_registers_i/depc_d [0]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_072_  (.A0(\i_ibex/csr_depc [10]),
    .A1(\i_ibex/cs_registers_i/depc_d [10]),
    .S(net921),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_073_  (.A0(\i_ibex/csr_depc [11]),
    .A1(\i_ibex/cs_registers_i/depc_d [11]),
    .S(net921),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_074_  (.A0(\i_ibex/csr_depc [12]),
    .A1(\i_ibex/cs_registers_i/depc_d [12]),
    .S(net921),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_075_  (.A0(\i_ibex/csr_depc [13]),
    .A1(\i_ibex/cs_registers_i/depc_d [13]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_076_  (.A0(\i_ibex/csr_depc [14]),
    .A1(\i_ibex/cs_registers_i/depc_d [14]),
    .S(net921),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_077_  (.A0(\i_ibex/csr_depc [15]),
    .A1(\i_ibex/cs_registers_i/depc_d [15]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_078_  (.A0(\i_ibex/csr_depc [16]),
    .A1(\i_ibex/cs_registers_i/depc_d [16]),
    .S(net923),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_079_  (.A0(\i_ibex/csr_depc [17]),
    .A1(\i_ibex/cs_registers_i/depc_d [17]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_080_  (.A0(\i_ibex/csr_depc [18]),
    .A1(\i_ibex/cs_registers_i/depc_d [18]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout861 (.A(net862),
    .X(net861),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_082_  (.A0(\i_ibex/csr_depc [19]),
    .A1(\i_ibex/cs_registers_i/depc_d [19]),
    .S(net923),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_083_  (.A0(\i_ibex/csr_depc [1]),
    .A1(\i_ibex/cs_registers_i/depc_d [1]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_084_  (.A0(\i_ibex/csr_depc [20]),
    .A1(\i_ibex/cs_registers_i/depc_d [20]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_085_  (.A0(\i_ibex/csr_depc [21]),
    .A1(\i_ibex/cs_registers_i/depc_d [21]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_086_  (.A0(\i_ibex/csr_depc [22]),
    .A1(\i_ibex/cs_registers_i/depc_d [22]),
    .S(net923),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_087_  (.A0(\i_ibex/csr_depc [23]),
    .A1(\i_ibex/cs_registers_i/depc_d [23]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_088_  (.A0(\i_ibex/csr_depc [24]),
    .A1(\i_ibex/cs_registers_i/depc_d [24]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_089_  (.A0(\i_ibex/csr_depc [25]),
    .A1(\i_ibex/cs_registers_i/depc_d [25]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_090_  (.A0(\i_ibex/csr_depc [26]),
    .A1(\i_ibex/cs_registers_i/depc_d [26]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_091_  (.A0(\i_ibex/csr_depc [27]),
    .A1(\i_ibex/cs_registers_i/depc_d [27]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout860 (.A(net394),
    .X(net860),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_093_  (.A0(\i_ibex/csr_depc [28]),
    .A1(\i_ibex/cs_registers_i/depc_d [28]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_094_  (.A0(\i_ibex/csr_depc [29]),
    .A1(\i_ibex/cs_registers_i/depc_d [29]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_095_  (.A0(\i_ibex/csr_depc [2]),
    .A1(\i_ibex/cs_registers_i/depc_d [2]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_096_  (.A0(\i_ibex/csr_depc [30]),
    .A1(\i_ibex/cs_registers_i/depc_d [30]),
    .S(net922),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_097_  (.A0(\i_ibex/csr_depc [31]),
    .A1(\i_ibex/cs_registers_i/depc_d [31]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_098_  (.A0(\i_ibex/csr_depc [3]),
    .A1(\i_ibex/cs_registers_i/depc_d [3]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_099_  (.A0(\i_ibex/csr_depc [4]),
    .A1(\i_ibex/cs_registers_i/depc_d [4]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_100_  (.A0(\i_ibex/csr_depc [5]),
    .A1(\i_ibex/cs_registers_i/depc_d [5]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_101_  (.A0(\i_ibex/csr_depc [6]),
    .A1(\i_ibex/cs_registers_i/depc_d [6]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_102_  (.A0(\i_ibex/csr_depc [7]),
    .A1(\i_ibex/cs_registers_i/depc_d [7]),
    .S(net920),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_103_  (.A0(\i_ibex/csr_depc [8]),
    .A1(\i_ibex/cs_registers_i/depc_d [8]),
    .S(net924),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_depc_csr/_104_  (.A0(\i_ibex/csr_depc [9]),
    .A1(\i_ibex/cs_registers_i/depc_d [9]),
    .S(net921),
    .X(\i_ibex/cs_registers_i/u_depc_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1440__66  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net66));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_76_clk_i_regs),
    .RESET_B(net1547),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_067_ ),
    .Q(\i_ibex/csr_depc [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[10]_reg  (.RESET_B(net1533),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_001_ ),
    .Q(\i_ibex/csr_depc [10]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_066_ ),
    .CLK(clknet_leaf_95_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[11]_reg  (.RESET_B(net1533),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_002_ ),
    .Q(\i_ibex/csr_depc [11]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_065_ ),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[12]_reg  (.RESET_B(net1568),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_003_ ),
    .Q(\i_ibex/csr_depc [12]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_064_ ),
    .CLK(clknet_leaf_80_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[13]_reg  (.RESET_B(net1593),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_004_ ),
    .Q(\i_ibex/csr_depc [13]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_063_ ),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[14]_reg  (.RESET_B(net1568),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_005_ ),
    .Q(\i_ibex/csr_depc [14]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_062_ ),
    .CLK(clknet_leaf_80_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_38_clk_i_regs),
    .RESET_B(net1593),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_061_ ),
    .Q(\i_ibex/csr_depc [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[16]_reg  (.RESET_B(net1626),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_007_ ),
    .Q(\i_ibex/csr_depc [16]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_060_ ),
    .CLK(clknet_leaf_139_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[17]_reg  (.RESET_B(net1633),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_008_ ),
    .Q(\i_ibex/csr_depc [17]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_059_ ),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[18]_reg  (.RESET_B(net1650),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_009_ ),
    .Q(\i_ibex/csr_depc [18]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_058_ ),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[19]_reg  (.RESET_B(net1654),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_010_ ),
    .Q(\i_ibex/csr_depc [19]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_057_ ),
    .CLK(clknet_leaf_139_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[1]_reg  (.RESET_B(net1572),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_011_ ),
    .Q(\i_ibex/csr_depc [1]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_056_ ),
    .CLK(clknet_leaf_75_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[20]_reg  (.RESET_B(net1625),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_012_ ),
    .Q(\i_ibex/csr_depc [20]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_055_ ),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[21]_reg  (.RESET_B(net1646),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_013_ ),
    .Q(\i_ibex/csr_depc [21]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_054_ ),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_28_clk_i_regs),
    .RESET_B(net1626),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_053_ ),
    .Q(\i_ibex/csr_depc [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_27_clk_i_regs),
    .RESET_B(net1646),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_052_ ),
    .Q(\i_ibex/csr_depc [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_28_clk_i_regs),
    .RESET_B(net1646),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_051_ ),
    .Q(\i_ibex/csr_depc [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_29_clk_i_regs),
    .RESET_B(net1648),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_050_ ),
    .Q(\i_ibex/csr_depc [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_29_clk_i_regs),
    .RESET_B(net1648),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_049_ ),
    .Q(\i_ibex/csr_depc [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_37_clk_i_regs),
    .RESET_B(net1592),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_048_ ),
    .Q(\i_ibex/csr_depc [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[28]_reg  (.RESET_B(net1596),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_020_ ),
    .Q(\i_ibex/csr_depc [28]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_047_ ),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_40_clk_i_regs),
    .RESET_B(net1605),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_046_ ),
    .Q(\i_ibex/csr_depc [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[2]_reg  (.RESET_B(net1570),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_022_ ),
    .Q(\i_ibex/csr_depc [2]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_045_ ),
    .CLK(clknet_leaf_78_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[30]_reg  (.RESET_B(net1646),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_023_ ),
    .Q(\i_ibex/csr_depc [30]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_044_ ),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[31]_reg  (.RESET_B(net1596),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_024_ ),
    .Q(\i_ibex/csr_depc [31]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_043_ ),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[3]_reg  (.RESET_B(net1570),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_025_ ),
    .Q(\i_ibex/csr_depc [3]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_042_ ),
    .CLK(clknet_leaf_78_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[4]_reg  (.RESET_B(net1572),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_026_ ),
    .Q(\i_ibex/csr_depc [4]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_041_ ),
    .CLK(clknet_leaf_75_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[5]_reg  (.RESET_B(net1569),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_027_ ),
    .Q(\i_ibex/csr_depc [5]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_040_ ),
    .CLK(clknet_leaf_81_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[6]_reg  (.RESET_B(net1569),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_028_ ),
    .Q(\i_ibex/csr_depc [6]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_039_ ),
    .CLK(clknet_leaf_81_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[7]_reg  (.RESET_B(net1569),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_029_ ),
    .Q(\i_ibex/csr_depc [7]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_038_ ),
    .CLK(clknet_leaf_81_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[8]_reg  (.RESET_B(net1604),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_030_ ),
    .Q(\i_ibex/csr_depc [8]),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_037_ ),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_depc_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1533),
    .D(\i_ibex/cs_registers_i/u_depc_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_depc_csr/_036_ ),
    .Q(\i_ibex/csr_depc [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout859 (.A(net860),
    .X(net859),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout858 (.A(net859),
    .X(net858),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_071_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [0]),
    .A1(net974),
    .S(net860),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_072_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [10]),
    .A1(net935),
    .S(net859),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_073_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [11]),
    .A1(net937),
    .S(net860),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_074_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [12]),
    .A1(net939),
    .S(net860),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_075_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [13]),
    .A1(net958),
    .S(net859),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_076_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [14]),
    .A1(net940),
    .S(net860),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_077_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [15]),
    .A1(net959),
    .S(net859),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_078_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [16]),
    .A1(net941),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_079_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [17]),
    .A1(net944),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_080_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [18]),
    .A1(net945),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout857 (.A(net858),
    .X(net857),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_082_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [19]),
    .A1(net947),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_083_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [1]),
    .A1(net972),
    .S(net860),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_084_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [20]),
    .A1(net427),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_085_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [21]),
    .A1(net962),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_086_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [22]),
    .A1(net413),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_087_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [23]),
    .A1(net415),
    .S(net857),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_088_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [24]),
    .A1(net927),
    .S(net858),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_089_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [25]),
    .A1(net417),
    .S(net858),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_090_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [26]),
    .A1(net929),
    .S(net858),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_091_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [27]),
    .A1(net424),
    .S(net892),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(\i_ibex/cs_registers_i/dcsr_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_093_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [28]),
    .A1(net418),
    .S(net892),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_094_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [29]),
    .A1(net420),
    .S(net892),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_095_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [2]),
    .A1(net950),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_096_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [30]),
    .A1(net964),
    .S(net892),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_097_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [31]),
    .A1(net423),
    .S(net892),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_098_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [3]),
    .A1(net951),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_099_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [4]),
    .A1(net954),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_100_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [5]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_101_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [6]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_102_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [7]),
    .A1(net955),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_103_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [8]),
    .A1(net931),
    .S(net892),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch0_csr/_104_  (.A0(\i_ibex/cs_registers_i/dscratch0_q [9]),
    .A1(net933),
    .S(net891),
    .X(\i_ibex/cs_registers_i/u_dscratch0_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1431__65  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net65));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_69_clk_i_regs),
    .RESET_B(net1540),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_067_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1603),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_001_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1602),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_065_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1602),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_064_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_52_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_004_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_063_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1608),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_53_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_6_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_6_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_6_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_71_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_056_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1639),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1640),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_24_clk_i_regs),
    .RESET_B(net1617),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_053_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1616),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_052_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1620),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_050_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_049_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1600),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_7_clk_i_regs),
    .RESET_B(net1616),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_047_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_46_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_046_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1538),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_045_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[30]_reg  (.CLK(clknet_leaf_6_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_044_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_19_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_043_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_69_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_041_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1535),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_040_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_039_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_038_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_037_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch0_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_61_clk_i_regs),
    .RESET_B(net1603),
    .D(\i_ibex/cs_registers_i/u_dscratch0_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch0_csr/_036_ ),
    .Q(\i_ibex/cs_registers_i/dscratch0_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(net856),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net855),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_071_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [0]),
    .A1(net974),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_072_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [10]),
    .A1(net935),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_073_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [11]),
    .A1(net937),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_074_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [12]),
    .A1(net939),
    .S(net906),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_075_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [13]),
    .A1(net958),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_076_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [14]),
    .A1(net940),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_077_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [15]),
    .A1(net959),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_078_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [16]),
    .A1(net941),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_079_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [17]),
    .A1(net944),
    .S(net904),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_080_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [18]),
    .A1(net945),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(\i_ibex/cs_registers_i/dcsr_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_082_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [19]),
    .A1(net947),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_083_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [1]),
    .A1(net972),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_084_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [20]),
    .A1(net427),
    .S(net904),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_085_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [21]),
    .A1(net962),
    .S(net904),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_086_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [22]),
    .A1(net413),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_087_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [23]),
    .A1(net415),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_088_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [24]),
    .A1(net927),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_089_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [25]),
    .A1(net417),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_090_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [26]),
    .A1(net929),
    .S(net904),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_091_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [27]),
    .A1(net424),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_093_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [28]),
    .A1(net419),
    .S(net903),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_094_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [29]),
    .A1(net420),
    .S(net905),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_095_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [2]),
    .A1(net950),
    .S(net906),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_096_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [30]),
    .A1(net964),
    .S(net904),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_097_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [31]),
    .A1(net423),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_098_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [3]),
    .A1(net951),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_099_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [4]),
    .A1(net954),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_100_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [5]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_101_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [6]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_102_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [7]),
    .A1(net955),
    .S(net901),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_103_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [8]),
    .A1(net931),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_dscratch1_csr/_104_  (.A0(\i_ibex/cs_registers_i/dscratch1_q [9]),
    .A1(net933),
    .S(net902),
    .X(\i_ibex/cs_registers_i/u_dscratch1_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1430__64  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net64));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_69_clk_i_regs),
    .RESET_B(net1540),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_067_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1603),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_001_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_61_clk_i_regs),
    .RESET_B(net1603),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_065_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1603),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_064_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1636),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_004_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_063_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1608),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1636),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_14_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_5_clk_i_regs),
    .RESET_B(net1645),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_19_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1649),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_056_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_3_clk_i_regs),
    .RESET_B(net1640),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_5_clk_i_regs),
    .RESET_B(net1645),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_19_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_053_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_052_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_18_clk_i_regs),
    .RESET_B(net1620),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_18_clk_i_regs),
    .RESET_B(net1620),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_050_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_19_clk_i_regs),
    .RESET_B(net1620),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_049_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1589),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_18_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_047_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_046_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1608),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_045_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[30]_reg  (.CLK(clknet_leaf_6_clk_i_regs),
    .RESET_B(net1645),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_044_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_043_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_041_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_67_clk_i_regs),
    .RESET_B(net1540),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_040_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1535),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_039_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1540),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_038_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1600),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_037_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_dscratch1_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_61_clk_i_regs),
    .RESET_B(net1600),
    .D(\i_ibex/cs_registers_i/u_dscratch1_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_dscratch1_csr/_036_ ),
    .Q(\i_ibex/cs_registers_i/dscratch1_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(net853),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_17_  (.A0(\i_ibex/cs_registers_i/mcause_q [0]),
    .A1(\i_ibex/cs_registers_i/mcause_d [0]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_00_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_18_  (.A0(\i_ibex/cs_registers_i/mcause_q [1]),
    .A1(\i_ibex/cs_registers_i/mcause_d [1]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_01_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_19_  (.A0(\i_ibex/cs_registers_i/mcause_q [2]),
    .A1(\i_ibex/cs_registers_i/mcause_d [2]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_02_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_20_  (.A0(\i_ibex/cs_registers_i/mcause_q [3]),
    .A1(\i_ibex/cs_registers_i/mcause_d [3]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_03_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_21_  (.A0(\i_ibex/cs_registers_i/mcause_q [4]),
    .A1(\i_ibex/cs_registers_i/mcause_d [4]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_04_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_22_  (.A0(\i_ibex/cs_registers_i/mcause_q [5]),
    .A1(\i_ibex/cs_registers_i/mcause_d [5]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_05_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mcause_csr/_23_  (.A0(\i_ibex/cs_registers_i/mcause_q [6]),
    .A1(\i_ibex/cs_registers_i/mcause_d [6]),
    .S(\i_ibex/cs_registers_i/mcause_en ),
    .X(\i_ibex/cs_registers_i/u_mcause_csr/_06_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1417__63  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net63));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_76_clk_i_regs),
    .RESET_B(net1547),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_00_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_14_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_72_clk_i_regs),
    .RESET_B(net1571),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_01_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_13_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_72_clk_i_regs),
    .RESET_B(net1571),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_02_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_12_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_72_clk_i_regs),
    .RESET_B(net1543),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_03_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_11_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_73_clk_i_regs),
    .RESET_B(net1548),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_04_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_10_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_76_clk_i_regs),
    .RESET_B(net1547),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_05_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_09_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mcause_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_78_clk_i_regs),
    .RESET_B(net1546),
    .D(\i_ibex/cs_registers_i/u_mcause_csr/_06_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mcause_csr/_08_ ),
    .Q(\i_ibex/cs_registers_i/mcause_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout850 (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_088_ ),
    .X(net850),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(net850),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_071_  (.A0(\i_ibex/csr_mepc [0]),
    .A1(\i_ibex/cs_registers_i/mepc_d [0]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_072_  (.A0(\i_ibex/csr_mepc [10]),
    .A1(\i_ibex/cs_registers_i/mepc_d [10]),
    .S(net881),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_073_  (.A0(\i_ibex/csr_mepc [11]),
    .A1(\i_ibex/cs_registers_i/mepc_d [11]),
    .S(net881),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_074_  (.A0(\i_ibex/csr_mepc [12]),
    .A1(\i_ibex/cs_registers_i/mepc_d [12]),
    .S(net881),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_075_  (.A0(\i_ibex/csr_mepc [13]),
    .A1(\i_ibex/cs_registers_i/mepc_d [13]),
    .S(net884),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_076_  (.A0(\i_ibex/csr_mepc [14]),
    .A1(\i_ibex/cs_registers_i/mepc_d [14]),
    .S(net881),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_077_  (.A0(\i_ibex/csr_mepc [15]),
    .A1(\i_ibex/cs_registers_i/mepc_d [15]),
    .S(net884),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_078_  (.A0(\i_ibex/csr_mepc [16]),
    .A1(\i_ibex/cs_registers_i/mepc_d [16]),
    .S(net883),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_079_  (.A0(\i_ibex/csr_mepc [17]),
    .A1(\i_ibex/cs_registers_i/mepc_d [17]),
    .S(net883),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_080_  (.A0(\i_ibex/csr_mepc [18]),
    .A1(\i_ibex/cs_registers_i/mepc_d [18]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout848 (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_173_ ),
    .X(net848),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_082_  (.A0(\i_ibex/csr_mepc [19]),
    .A1(\i_ibex/cs_registers_i/mepc_d [19]),
    .S(net883),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_083_  (.A0(\i_ibex/csr_mepc [1]),
    .A1(\i_ibex/cs_registers_i/mepc_d [1]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_084_  (.A0(\i_ibex/csr_mepc [20]),
    .A1(\i_ibex/cs_registers_i/mepc_d [20]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_085_  (.A0(\i_ibex/csr_mepc [21]),
    .A1(\i_ibex/cs_registers_i/mepc_d [21]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_086_  (.A0(\i_ibex/csr_mepc [22]),
    .A1(\i_ibex/cs_registers_i/mepc_d [22]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_087_  (.A0(\i_ibex/csr_mepc [23]),
    .A1(\i_ibex/cs_registers_i/mepc_d [23]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_088_  (.A0(\i_ibex/csr_mepc [24]),
    .A1(\i_ibex/cs_registers_i/mepc_d [24]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_089_  (.A0(\i_ibex/csr_mepc [25]),
    .A1(\i_ibex/cs_registers_i/mepc_d [25]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_090_  (.A0(\i_ibex/csr_mepc [26]),
    .A1(\i_ibex/cs_registers_i/mepc_d [26]),
    .S(net882),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_091_  (.A0(\i_ibex/csr_mepc [27]),
    .A1(\i_ibex/cs_registers_i/mepc_d [27]),
    .S(net884),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout847 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0236_ ),
    .X(net847),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_093_  (.A0(\i_ibex/csr_mepc [28]),
    .A1(\i_ibex/cs_registers_i/mepc_d [28]),
    .S(net884),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_094_  (.A0(\i_ibex/csr_mepc [29]),
    .A1(\i_ibex/cs_registers_i/mepc_d [29]),
    .S(net884),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_095_  (.A0(\i_ibex/csr_mepc [2]),
    .A1(\i_ibex/cs_registers_i/mepc_d [2]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_096_  (.A0(\i_ibex/csr_mepc [30]),
    .A1(\i_ibex/cs_registers_i/mepc_d [30]),
    .S(net883),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_097_  (.A0(\i_ibex/csr_mepc [31]),
    .A1(\i_ibex/cs_registers_i/mepc_d [31]),
    .S(net883),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_098_  (.A0(\i_ibex/csr_mepc [3]),
    .A1(\i_ibex/cs_registers_i/mepc_d [3]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_099_  (.A0(\i_ibex/csr_mepc [4]),
    .A1(\i_ibex/cs_registers_i/mepc_d [4]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_100_  (.A0(\i_ibex/csr_mepc [5]),
    .A1(\i_ibex/cs_registers_i/mepc_d [5]),
    .S(net881),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_101_  (.A0(\i_ibex/csr_mepc [6]),
    .A1(\i_ibex/cs_registers_i/mepc_d [6]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_102_  (.A0(\i_ibex/csr_mepc [7]),
    .A1(\i_ibex/cs_registers_i/mepc_d [7]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_103_  (.A0(\i_ibex/csr_mepc [8]),
    .A1(\i_ibex/cs_registers_i/mepc_d [8]),
    .S(net880),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mepc_csr/_104_  (.A0(\i_ibex/csr_mepc [9]),
    .A1(\i_ibex/cs_registers_i/mepc_d [9]),
    .S(net881),
    .X(\i_ibex/cs_registers_i/u_mepc_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1416__62  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net62));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_73_clk_i_regs),
    .RESET_B(net1543),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_067_ ),
    .Q(\i_ibex/csr_mepc [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[10]_reg  (.RESET_B(net1533),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_001_ ),
    .Q(\i_ibex/csr_mepc [10]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_066_ ),
    .CLK(clknet_leaf_94_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[11]_reg  (.RESET_B(net1550),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_002_ ),
    .Q(\i_ibex/csr_mepc [11]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_065_ ),
    .CLK(clknet_leaf_94_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[12]_reg  (.RESET_B(net1568),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_003_ ),
    .Q(\i_ibex/csr_mepc [12]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_064_ ),
    .CLK(clknet_leaf_82_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[13]_reg  (.RESET_B(net1593),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_004_ ),
    .Q(\i_ibex/csr_mepc [13]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_063_ ),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[14]_reg  (.RESET_B(net1568),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_005_ ),
    .Q(\i_ibex/csr_mepc [14]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_062_ ),
    .CLK(clknet_leaf_93_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[15]_reg  (.RESET_B(net1593),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_006_ ),
    .Q(\i_ibex/csr_mepc [15]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_061_ ),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_31_clk_i_regs),
    .RESET_B(net1633),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_060_ ),
    .Q(\i_ibex/csr_mepc [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[17]_reg  (.RESET_B(net1655),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_008_ ),
    .Q(\i_ibex/csr_mepc [17]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_059_ ),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[18]_reg  (.RESET_B(net1654),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_009_ ),
    .Q(\i_ibex/csr_mepc [18]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_058_ ),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[19]_reg  (.RESET_B(net1655),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_010_ ),
    .Q(\i_ibex/csr_mepc [19]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_057_ ),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[1]_reg  (.RESET_B(net1571),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_011_ ),
    .Q(\i_ibex/csr_mepc [1]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_056_ ),
    .CLK(clknet_leaf_73_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[20]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_012_ ),
    .Q(\i_ibex/csr_mepc [20]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_055_ ),
    .CLK(clknet_leaf_139_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[21]_reg  (.RESET_B(net1652),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_013_ ),
    .Q(\i_ibex/csr_mepc [21]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_054_ ),
    .CLK(clknet_leaf_138_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[22]_reg  (.RESET_B(net1626),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_014_ ),
    .Q(\i_ibex/csr_mepc [22]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_053_ ),
    .CLK(clknet_leaf_137_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[23]_reg  (.RESET_B(net1626),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_015_ ),
    .Q(\i_ibex/csr_mepc [23]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_052_ ),
    .CLK(clknet_leaf_137_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[24]_reg  (.RESET_B(net1653),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_016_ ),
    .Q(\i_ibex/csr_mepc [24]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_051_ ),
    .CLK(clknet_leaf_139_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[25]_reg  (.RESET_B(net1654),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_017_ ),
    .Q(\i_ibex/csr_mepc [25]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_050_ ),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[26]_reg  (.RESET_B(net1654),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_018_ ),
    .Q(\i_ibex/csr_mepc [26]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_049_ ),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[27]_reg  (.RESET_B(net1592),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_019_ ),
    .Q(\i_ibex/csr_mepc [27]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_048_ ),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_34_clk_i_regs),
    .RESET_B(net1592),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_047_ ),
    .Q(\i_ibex/csr_mepc [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_41_clk_i_regs),
    .RESET_B(net1605),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_046_ ),
    .Q(\i_ibex/csr_mepc [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[2]_reg  (.RESET_B(net1572),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_022_ ),
    .Q(\i_ibex/csr_mepc [2]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_045_ ),
    .CLK(clknet_leaf_73_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[30]_reg  (.RESET_B(net1655),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_023_ ),
    .Q(\i_ibex/csr_mepc [30]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_044_ ),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[31]_reg  (.RESET_B(net1633),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_024_ ),
    .Q(\i_ibex/csr_mepc [31]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_043_ ),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[3]_reg  (.RESET_B(net1574),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_025_ ),
    .Q(\i_ibex/csr_mepc [3]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_042_ ),
    .CLK(clknet_leaf_74_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[4]_reg  (.RESET_B(net1571),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_026_ ),
    .Q(\i_ibex/csr_mepc [4]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_041_ ),
    .CLK(clknet_leaf_74_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[5]_reg  (.RESET_B(net1573),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_027_ ),
    .Q(\i_ibex/csr_mepc [5]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_040_ ),
    .CLK(clknet_leaf_84_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[6]_reg  (.RESET_B(net1573),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_028_ ),
    .Q(\i_ibex/csr_mepc [6]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_039_ ),
    .CLK(clknet_leaf_84_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[7]_reg  (.RESET_B(net1574),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_029_ ),
    .Q(\i_ibex/csr_mepc [7]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_038_ ),
    .CLK(clknet_leaf_85_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[8]_reg  (.RESET_B(net1547),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_030_ ),
    .Q(\i_ibex/csr_mepc [8]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_037_ ),
    .CLK(clknet_leaf_75_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mepc_csr/rd_data_o[9]_reg  (.RESET_B(net1546),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mepc_csr/_031_ ),
    .Q(\i_ibex/csr_mepc [9]),
    .Q_N(\i_ibex/cs_registers_i/u_mepc_csr/_036_ ),
    .CLK(clknet_leaf_94_clk_i_regs));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0236_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout845 (.X(net845),
    .A(\i_ibex/if_stage_i/_340_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_43_  (.A0(\i_ibex/cs_registers_i/mie_q [0]),
    .A1(net941),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_00_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_44_  (.A0(\i_ibex/cs_registers_i/mie_q [10]),
    .A1(net929),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_01_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_45_  (.A0(\i_ibex/cs_registers_i/mie_q [11]),
    .A1(net424),
    .S(net900),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_02_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_46_  (.A0(\i_ibex/cs_registers_i/mie_q [12]),
    .A1(net419),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_03_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_47_  (.A0(\i_ibex/cs_registers_i/mie_q [13]),
    .A1(net420),
    .S(net900),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_04_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_48_  (.A0(\i_ibex/cs_registers_i/mie_q [14]),
    .A1(net964),
    .S(net899),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_05_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_49_  (.A0(\i_ibex/cs_registers_i/mie_q [15]),
    .A1(net423),
    .S(net899),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_06_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_50_  (.A0(\i_ibex/cs_registers_i/mie_q [16]),
    .A1(net938),
    .S(net900),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_07_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_51_  (.A0(\i_ibex/cs_registers_i/mie_q [17]),
    .A1(net956),
    .S(net900),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_08_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_52_  (.A0(\i_ibex/cs_registers_i/mie_q [18]),
    .A1(net952),
    .S(net900),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_09_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_53_  (.A0(\i_ibex/cs_registers_i/mie_q [1]),
    .A1(net943),
    .S(net900),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_10_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_54_  (.A0(\i_ibex/cs_registers_i/mie_q [2]),
    .A1(net945),
    .S(net899),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_11_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_55_  (.A0(\i_ibex/cs_registers_i/mie_q [3]),
    .A1(net947),
    .S(net899),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_12_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_56_  (.A0(\i_ibex/cs_registers_i/mie_q [4]),
    .A1(net427),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_13_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_57_  (.A0(\i_ibex/cs_registers_i/mie_q [5]),
    .A1(net961),
    .S(net899),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_14_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_58_  (.A0(\i_ibex/cs_registers_i/mie_q [6]),
    .A1(net413),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_15_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_59_  (.A0(\i_ibex/cs_registers_i/mie_q [7]),
    .A1(net415),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_16_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_60_  (.A0(\i_ibex/cs_registers_i/mie_q [8]),
    .A1(net927),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_17_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mie_csr/_61_  (.A0(\i_ibex/cs_registers_i/mie_q [9]),
    .A1(net417),
    .S(net898),
    .X(\i_ibex/cs_registers_i/u_mie_csr/_18_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1409__61  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net61));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_00_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_39_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_24_clk_i_regs),
    .RESET_B(net1620),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_01_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_38_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1591),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_02_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_37_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_03_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_36_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_50_clk_i_regs),
    .RESET_B(net1599),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_04_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_35_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1622),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_05_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_34_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[15]_reg  (.RESET_B(net1589),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_06_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [15]),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_33_ ),
    .CLK(clknet_leaf_49_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_46_clk_i_regs),
    .RESET_B(net1604),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_07_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_32_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_45_clk_i_regs),
    .RESET_B(net1531),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_08_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_31_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_45_clk_i_regs),
    .RESET_B(net1531),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_09_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_30_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_47_clk_i_regs),
    .RESET_B(net1604),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_10_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_29_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_21_clk_i_regs),
    .RESET_B(net1622),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_11_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_28_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1621),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_12_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_27_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_20_clk_i_regs),
    .RESET_B(net1632),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_13_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_26_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1589),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_14_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_25_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_19_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_15_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_24_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_19_clk_i_regs),
    .RESET_B(net1620),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_16_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_23_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_24_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_17_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_22_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mie_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_24_clk_i_regs),
    .RESET_B(net1619),
    .D(\i_ibex/cs_registers_i/u_mie_csr/_18_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mie_csr/_21_ ),
    .Q(\i_ibex/cs_registers_i/mie_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(net845),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net844),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_071_  (.A0(\i_ibex/cs_registers_i/mscratch_q [0]),
    .A1(net974),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_072_  (.A0(\i_ibex/cs_registers_i/mscratch_q [10]),
    .A1(net935),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_073_  (.A0(\i_ibex/cs_registers_i/mscratch_q [11]),
    .A1(net938),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_074_  (.A0(\i_ibex/cs_registers_i/mscratch_q [12]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [12]),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_075_  (.A0(\i_ibex/cs_registers_i/mscratch_q [13]),
    .A1(net957),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_076_  (.A0(\i_ibex/cs_registers_i/mscratch_q [14]),
    .A1(net940),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_077_  (.A0(\i_ibex/cs_registers_i/mscratch_q [15]),
    .A1(net959),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_078_  (.A0(\i_ibex/cs_registers_i/mscratch_q [16]),
    .A1(net942),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_079_  (.A0(\i_ibex/cs_registers_i/mscratch_q [17]),
    .A1(net944),
    .S(net873),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_080_  (.A0(\i_ibex/cs_registers_i/mscratch_q [18]),
    .A1(net946),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(\i_ibex/if_stage_i/_340_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_082_  (.A0(\i_ibex/cs_registers_i/mscratch_q [19]),
    .A1(net948),
    .S(net873),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_083_  (.A0(\i_ibex/cs_registers_i/mscratch_q [1]),
    .A1(net972),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_084_  (.A0(\i_ibex/cs_registers_i/mscratch_q [20]),
    .A1(net427),
    .S(net874),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_085_  (.A0(\i_ibex/cs_registers_i/mscratch_q [21]),
    .A1(net962),
    .S(net873),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_086_  (.A0(\i_ibex/cs_registers_i/mscratch_q [22]),
    .A1(net413),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_087_  (.A0(\i_ibex/cs_registers_i/mscratch_q [23]),
    .A1(net415),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_088_  (.A0(\i_ibex/cs_registers_i/mscratch_q [24]),
    .A1(net928),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_089_  (.A0(\i_ibex/cs_registers_i/mscratch_q [25]),
    .A1(net417),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_090_  (.A0(\i_ibex/cs_registers_i/mscratch_q [26]),
    .A1(net930),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_091_  (.A0(\i_ibex/cs_registers_i/mscratch_q [27]),
    .A1(net425),
    .S(net874),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(net842),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_093_  (.A0(\i_ibex/cs_registers_i/mscratch_q [28]),
    .A1(net419),
    .S(net873),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_094_  (.A0(\i_ibex/cs_registers_i/mscratch_q [29]),
    .A1(net421),
    .S(net874),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_095_  (.A0(\i_ibex/cs_registers_i/mscratch_q [2]),
    .A1(net949),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_096_  (.A0(\i_ibex/cs_registers_i/mscratch_q [30]),
    .A1(net964),
    .S(net872),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_097_  (.A0(\i_ibex/cs_registers_i/mscratch_q [31]),
    .A1(net423),
    .S(net871),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_098_  (.A0(\i_ibex/cs_registers_i/mscratch_q [3]),
    .A1(net951),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_099_  (.A0(\i_ibex/cs_registers_i/mscratch_q [4]),
    .A1(net954),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_100_  (.A0(\i_ibex/cs_registers_i/mscratch_q [5]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [5]),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_101_  (.A0(\i_ibex/cs_registers_i/mscratch_q [6]),
    .A1(\i_ibex/cs_registers_i/csr_wdata_int [6]),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_102_  (.A0(\i_ibex/cs_registers_i/mscratch_q [7]),
    .A1(net956),
    .S(net875),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_103_  (.A0(\i_ibex/cs_registers_i/mscratch_q [8]),
    .A1(net932),
    .S(net870),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mscratch_csr/_104_  (.A0(\i_ibex/cs_registers_i/mscratch_q [9]),
    .A1(net934),
    .S(net875),
    .X(\i_ibex/cs_registers_i/u_mscratch_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1408__60  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net60));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_067_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1529),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_001_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_79_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_065_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_77_clk_i_regs),
    .RESET_B(net1538),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_064_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_61_clk_i_regs),
    .RESET_B(net1529),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_004_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_063_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_61_clk_i_regs),
    .RESET_B(net1552),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_48_clk_i_regs),
    .RESET_B(net1595),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_76_clk_i_regs),
    .RESET_B(net1542),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_056_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_48_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_48_clk_i_regs),
    .RESET_B(net1632),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1630),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_053_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_23_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_052_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_23_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_23_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_050_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_23_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_049_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_49_clk_i_regs),
    .RESET_B(net1589),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_22_clk_i_regs),
    .RESET_B(net1631),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_047_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_47_clk_i_regs),
    .RESET_B(net1604),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_046_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1539),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_045_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[30]_reg  (.CLK(clknet_leaf_23_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_044_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_62_clk_i_regs),
    .RESET_B(net1538),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_043_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_77_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_77_clk_i_regs),
    .RESET_B(net1541),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_041_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_78_clk_i_regs),
    .RESET_B(net1546),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_040_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1538),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_039_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_45_clk_i_regs),
    .RESET_B(net1532),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_038_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_78_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_037_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mscratch_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1532),
    .D(\i_ibex/cs_registers_i/u_mscratch_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mscratch_csr/_036_ ),
    .Q(\i_ibex/cs_registers_i/mscratch_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout840 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_176_ ),
    .X(net840),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_17_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [0]),
    .A1(\i_ibex/cs_registers_i/mcause_q [0]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_00_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_18_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [1]),
    .A1(\i_ibex/cs_registers_i/mcause_q [1]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_01_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_19_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [2]),
    .A1(\i_ibex/cs_registers_i/mcause_q [2]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_02_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_20_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [3]),
    .A1(\i_ibex/cs_registers_i/mcause_q [3]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_03_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_21_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [4]),
    .A1(\i_ibex/cs_registers_i/mcause_q [4]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_04_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_22_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [5]),
    .A1(\i_ibex/cs_registers_i/mcause_q [5]),
    .S(net1045),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_05_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/_23_  (.A0(\i_ibex/cs_registers_i/mstack_cause_q [6]),
    .A1(\i_ibex/cs_registers_i/mcause_q [6]),
    .S(net1046),
    .X(\i_ibex/cs_registers_i/u_mstack_cause_csr/_06_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1404__59  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net59));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_76_clk_i_regs),
    .RESET_B(net1572),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_00_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_14_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_72_clk_i_regs),
    .RESET_B(net1571),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_01_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_13_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_71_clk_i_regs),
    .RESET_B(net1572),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_02_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_12_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_73_clk_i_regs),
    .RESET_B(net1543),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_03_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_11_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_73_clk_i_regs),
    .RESET_B(net1548),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_04_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_10_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_75_clk_i_regs),
    .RESET_B(net1572),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_05_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_09_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_cause_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_81_clk_i_regs),
    .RESET_B(net1550),
    .D(\i_ibex/cs_registers_i/u_mstack_cause_csr/_06_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_cause_csr/_08_ ),
    .Q(\i_ibex/cs_registers_i/mstack_cause_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_csr/_08_  (.A0(\i_ibex/cs_registers_i/mstack_q [0]),
    .A1(\i_ibex/cs_registers_i/mstatus_q [2]),
    .S(net1045),
    .X(\i_ibex/cs_registers_i/u_mstack_csr/_01_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_csr/_09_  (.A0(\i_ibex/cs_registers_i/mstack_q [1]),
    .A1(\i_ibex/cs_registers_i/mstatus_q [3]),
    .S(net1045),
    .X(\i_ibex/cs_registers_i/u_mstack_csr/_02_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_mstack_csr/_10_  (.A(\i_ibex/cs_registers_i/u_mstack_csr/_00_ ),
    .B(net1056),
    .Y(\i_ibex/cs_registers_i/u_mstack_csr/_04_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_mstack_csr/_11_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mstatus_q [4]),
    .A2(net1056),
    .Y(\i_ibex/cs_registers_i/u_mstack_csr/_03_ ),
    .B1(\i_ibex/cs_registers_i/u_mstack_csr/_04_ ));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1403__58  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net58));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_74_clk_i_regs),
    .RESET_B(net1547),
    .D(\i_ibex/cs_registers_i/u_mstack_csr/_01_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_csr/_06_ ),
    .Q(\i_ibex/cs_registers_i/mstack_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_85_clk_i_regs),
    .RESET_B(net1549),
    .D(\i_ibex/cs_registers_i/u_mstack_csr/_02_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_csr/_05_ ),
    .Q(\i_ibex/cs_registers_i/mstack_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_85_clk_i_regs),
    .RESET_B(net1573),
    .D(\i_ibex/cs_registers_i/u_mstack_csr/_03_ ),
    .Q_N(\i_ibex/cs_registers_i/mstack_q [2]),
    .Q(\i_ibex/cs_registers_i/u_mstack_csr/_00_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout839 (.X(net839),
    .A(net840),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout838 (.X(net838),
    .A(net839),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_071_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [0]),
    .A1(\i_ibex/csr_mepc [0]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_072_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [10]),
    .A1(\i_ibex/csr_mepc [10]),
    .S(net1046),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_073_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [11]),
    .A1(\i_ibex/csr_mepc [11]),
    .S(net1046),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_074_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [12]),
    .A1(\i_ibex/csr_mepc [12]),
    .S(net1046),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_075_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [13]),
    .A1(\i_ibex/csr_mepc [13]),
    .S(net1049),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_076_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [14]),
    .A1(\i_ibex/csr_mepc [14]),
    .S(net1046),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_077_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [15]),
    .A1(\i_ibex/csr_mepc [15]),
    .S(net1049),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_078_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [16]),
    .A1(\i_ibex/csr_mepc [16]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_079_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [17]),
    .A1(\i_ibex/csr_mepc [17]),
    .S(net1048),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_080_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [18]),
    .A1(\i_ibex/csr_mepc [18]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout837 (.X(net837),
    .A(net382),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_082_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [19]),
    .A1(\i_ibex/csr_mepc [19]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_083_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [1]),
    .A1(\i_ibex/csr_mepc [1]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_084_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [20]),
    .A1(\i_ibex/csr_mepc [20]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_085_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [21]),
    .A1(\i_ibex/csr_mepc [21]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_086_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [22]),
    .A1(\i_ibex/csr_mepc [22]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_087_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [23]),
    .A1(\i_ibex/csr_mepc [23]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_088_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [24]),
    .A1(\i_ibex/csr_mepc [24]),
    .S(net1047),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_089_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [25]),
    .A1(\i_ibex/csr_mepc [25]),
    .S(net1048),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_090_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [26]),
    .A1(\i_ibex/csr_mepc [26]),
    .S(net1048),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_091_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [27]),
    .A1(\i_ibex/csr_mepc [27]),
    .S(net1049),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout836 (.X(net836),
    .A(net837),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_093_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [28]),
    .A1(\i_ibex/csr_mepc [28]),
    .S(net1049),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_094_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [29]),
    .A1(\i_ibex/csr_mepc [29]),
    .S(net1049),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_095_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [2]),
    .A1(\i_ibex/csr_mepc [2]),
    .S(net1044),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_096_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [30]),
    .A1(\i_ibex/csr_mepc [30]),
    .S(net1048),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_097_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [31]),
    .A1(\i_ibex/csr_mepc [31]),
    .S(net1048),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_098_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [3]),
    .A1(\i_ibex/csr_mepc [3]),
    .S(net1044),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_099_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [4]),
    .A1(\i_ibex/csr_mepc [4]),
    .S(net1044),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_100_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [5]),
    .A1(\i_ibex/csr_mepc [5]),
    .S(net1045),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_101_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [6]),
    .A1(\i_ibex/csr_mepc [6]),
    .S(net1045),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_102_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [7]),
    .A1(\i_ibex/csr_mepc [7]),
    .S(net1044),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_103_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [8]),
    .A1(\i_ibex/csr_mepc [8]),
    .S(net1043),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/_104_  (.A0(\i_ibex/cs_registers_i/mstack_epc_q [9]),
    .A1(\i_ibex/csr_mepc [9]),
    .S(net1046),
    .X(\i_ibex/cs_registers_i/u_mstack_epc_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1396__57  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net57));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_72_clk_i_regs),
    .RESET_B(net1543),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_067_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_93_clk_i_regs),
    .RESET_B(net1546),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_001_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_93_clk_i_regs),
    .RESET_B(net1550),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_065_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_93_clk_i_regs),
    .RESET_B(net1568),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_064_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_37_clk_i_regs),
    .RESET_B(net1593),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_004_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_063_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_93_clk_i_regs),
    .RESET_B(net1568),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_37_clk_i_regs),
    .RESET_B(net1593),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_29_clk_i_regs),
    .RESET_B(net1626),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_30_clk_i_regs),
    .RESET_B(net1654),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_137_clk_i_regs),
    .RESET_B(net1654),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_29_clk_i_regs),
    .RESET_B(net1654),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_73_clk_i_regs),
    .RESET_B(net1571),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_056_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_138_clk_i_regs),
    .RESET_B(net1653),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_138_clk_i_regs),
    .RESET_B(net1652),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_137_clk_i_regs),
    .RESET_B(net1626),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_053_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_138_clk_i_regs),
    .RESET_B(net1652),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_052_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_139_clk_i_regs),
    .RESET_B(net1653),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_137_clk_i_regs),
    .RESET_B(net1655),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_050_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_30_clk_i_regs),
    .RESET_B(net1654),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_049_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_34_clk_i_regs),
    .RESET_B(net1592),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_34_clk_i_regs),
    .RESET_B(net1592),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_047_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_37_clk_i_regs),
    .RESET_B(net1593),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_046_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_73_clk_i_regs),
    .RESET_B(net1571),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_045_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[30]_reg  (.CLK(clknet_leaf_137_clk_i_regs),
    .RESET_B(net1655),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_044_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_31_clk_i_regs),
    .RESET_B(net1634),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_043_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_74_clk_i_regs),
    .RESET_B(net1548),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_74_clk_i_regs),
    .RESET_B(net1571),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_041_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_81_clk_i_regs),
    .RESET_B(net1569),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_040_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_84_clk_i_regs),
    .RESET_B(net1573),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_039_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_74_clk_i_regs),
    .RESET_B(net1572),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_038_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_75_clk_i_regs),
    .RESET_B(net1548),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_037_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mstack_epc_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_94_clk_i_regs),
    .RESET_B(net1546),
    .D(\i_ibex/cs_registers_i/u_mstack_epc_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mstack_epc_csr/_036_ ),
    .Q(\i_ibex/cs_registers_i/mstack_epc_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout835 (.X(net835),
    .A(net836),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstatus_csr/_17_  (.A0(\i_ibex/csr_mstatus_tw ),
    .A1(\i_ibex/cs_registers_i/mstatus_d [0]),
    .S(\i_ibex/cs_registers_i/mstatus_en ),
    .X(\i_ibex/cs_registers_i/u_mstatus_csr/_02_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstatus_csr/_18_  (.A0(\i_ibex/cs_registers_i/mstatus_q [1]),
    .A1(\i_ibex/cs_registers_i/mstatus_d [1]),
    .S(\i_ibex/cs_registers_i/mstatus_en ),
    .X(\i_ibex/cs_registers_i/u_mstatus_csr/_03_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_mstatus_csr/_19_  (.A(\i_ibex/cs_registers_i/u_mstatus_csr/_00_ ),
    .B(\i_ibex/cs_registers_i/mstatus_en ),
    .Y(\i_ibex/cs_registers_i/u_mstatus_csr/_09_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_mstatus_csr/_20_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mstatus_d [2]),
    .A2(\i_ibex/cs_registers_i/mstatus_en ),
    .Y(\i_ibex/cs_registers_i/u_mstatus_csr/_04_ ),
    .B1(\i_ibex/cs_registers_i/u_mstatus_csr/_09_ ));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_mstatus_csr/_21_  (.A(\i_ibex/cs_registers_i/u_mstatus_csr/_01_ ),
    .B(\i_ibex/cs_registers_i/mstatus_en ),
    .Y(\i_ibex/cs_registers_i/u_mstatus_csr/_10_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_mstatus_csr/_22_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/cs_registers_i/mstatus_d [3]),
    .A2(\i_ibex/cs_registers_i/mstatus_en ),
    .Y(\i_ibex/cs_registers_i/u_mstatus_csr/_05_ ),
    .B1(\i_ibex/cs_registers_i/u_mstatus_csr/_10_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstatus_csr/_23_  (.A0(\i_ibex/cs_registers_i/mstatus_q [4]),
    .A1(\i_ibex/cs_registers_i/mstatus_d [4]),
    .S(\i_ibex/cs_registers_i/mstatus_en ),
    .X(\i_ibex/cs_registers_i/u_mstatus_csr/_06_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mstatus_csr/_24_  (.A0(\i_ibex/csr_mstatus_mie ),
    .A1(\i_ibex/cs_registers_i/mstatus_d [5]),
    .S(\i_ibex/cs_registers_i/mstatus_en ),
    .X(\i_ibex/cs_registers_i/u_mstatus_csr/_07_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1395__56  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net56));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mstatus_csr/rd_data_o[0]_reg  (.RESET_B(net1573),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mstatus_csr/_02_ ),
    .Q(\i_ibex/csr_mstatus_tw ),
    .Q_N(\i_ibex/cs_registers_i/u_mstatus_csr/_14_ ),
    .CLK(clknet_leaf_84_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mstatus_csr/rd_data_o[1]_reg  (.RESET_B(net1547),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mstatus_csr/_03_ ),
    .Q(\i_ibex/cs_registers_i/mstatus_q [1]),
    .Q_N(\i_ibex/cs_registers_i/u_mstatus_csr/_13_ ),
    .CLK(clknet_leaf_75_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mstatus_csr/rd_data_o[2]_reg  (.RESET_B(net1547),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mstatus_csr/_04_ ),
    .Q(\i_ibex/cs_registers_i/u_mstatus_csr/_00_ ),
    .Q_N(\i_ibex/cs_registers_i/mstatus_q [2]),
    .CLK(clknet_leaf_74_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mstatus_csr/rd_data_o[3]_reg  (.RESET_B(net1548),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mstatus_csr/_05_ ),
    .Q(\i_ibex/cs_registers_i/u_mstatus_csr/_01_ ),
    .Q_N(\i_ibex/cs_registers_i/mstatus_q [3]),
    .CLK(clknet_leaf_74_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mstatus_csr/rd_data_o[4]_reg  (.RESET_B(net1573),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mstatus_csr/_06_ ),
    .Q(\i_ibex/cs_registers_i/mstatus_q [4]),
    .Q_N(\i_ibex/cs_registers_i/u_mstatus_csr/_12_ ),
    .CLK(clknet_leaf_85_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mstatus_csr/rd_data_o[5]_reg  (.RESET_B(net1574),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mstatus_csr/_07_ ),
    .Q(\i_ibex/csr_mstatus_mie ),
    .Q_N(\i_ibex/cs_registers_i/u_mstatus_csr/_11_ ),
    .CLK(clknet_leaf_85_clk_i_regs));
 sg13g2_buf_16 fanout834 (.X(net834),
    .A(net837),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout833 (.X(net833),
    .A(net834),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_071_  (.A0(\i_ibex/cs_registers_i/mtval_q [0]),
    .A1(\i_ibex/cs_registers_i/mtval_d [0]),
    .S(net869),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_072_  (.A0(\i_ibex/cs_registers_i/mtval_q [10]),
    .A1(\i_ibex/cs_registers_i/mtval_d [10]),
    .S(net865),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_073_  (.A0(\i_ibex/cs_registers_i/mtval_q [11]),
    .A1(\i_ibex/cs_registers_i/mtval_d [11]),
    .S(net866),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_074_  (.A0(\i_ibex/cs_registers_i/mtval_q [12]),
    .A1(\i_ibex/cs_registers_i/mtval_d [12]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_075_  (.A0(\i_ibex/cs_registers_i/mtval_q [13]),
    .A1(\i_ibex/cs_registers_i/mtval_d [13]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_076_  (.A0(\i_ibex/cs_registers_i/mtval_q [14]),
    .A1(\i_ibex/cs_registers_i/mtval_d [14]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_077_  (.A0(\i_ibex/cs_registers_i/mtval_q [15]),
    .A1(\i_ibex/cs_registers_i/mtval_d [15]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_078_  (.A0(\i_ibex/cs_registers_i/mtval_q [16]),
    .A1(\i_ibex/cs_registers_i/mtval_d [16]),
    .S(net868),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_079_  (.A0(\i_ibex/cs_registers_i/mtval_q [17]),
    .A1(\i_ibex/cs_registers_i/mtval_d [17]),
    .S(net869),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_080_  (.A0(\i_ibex/cs_registers_i/mtval_q [18]),
    .A1(\i_ibex/cs_registers_i/mtval_d [18]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout832 (.X(net832),
    .A(net834),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_082_  (.A0(\i_ibex/cs_registers_i/mtval_q [19]),
    .A1(\i_ibex/cs_registers_i/mtval_d [19]),
    .S(net868),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_083_  (.A0(\i_ibex/cs_registers_i/mtval_q [1]),
    .A1(\i_ibex/cs_registers_i/mtval_d [1]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_084_  (.A0(\i_ibex/cs_registers_i/mtval_q [20]),
    .A1(\i_ibex/cs_registers_i/mtval_d [20]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_085_  (.A0(\i_ibex/cs_registers_i/mtval_q [21]),
    .A1(\i_ibex/cs_registers_i/mtval_d [21]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_086_  (.A0(\i_ibex/cs_registers_i/mtval_q [22]),
    .A1(\i_ibex/cs_registers_i/mtval_d [22]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_087_  (.A0(\i_ibex/cs_registers_i/mtval_q [23]),
    .A1(\i_ibex/cs_registers_i/mtval_d [23]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_088_  (.A0(\i_ibex/cs_registers_i/mtval_q [24]),
    .A1(\i_ibex/cs_registers_i/mtval_d [24]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_089_  (.A0(\i_ibex/cs_registers_i/mtval_q [25]),
    .A1(\i_ibex/cs_registers_i/mtval_d [25]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_090_  (.A0(\i_ibex/cs_registers_i/mtval_q [26]),
    .A1(\i_ibex/cs_registers_i/mtval_d [26]),
    .S(net867),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_091_  (.A0(\i_ibex/cs_registers_i/mtval_q [27]),
    .A1(\i_ibex/cs_registers_i/mtval_d [27]),
    .S(net868),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout831 (.X(net831),
    .A(net832),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_093_  (.A0(\i_ibex/cs_registers_i/mtval_q [28]),
    .A1(\i_ibex/cs_registers_i/mtval_d [28]),
    .S(net869),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_094_  (.A0(\i_ibex/cs_registers_i/mtval_q [29]),
    .A1(\i_ibex/cs_registers_i/mtval_d [29]),
    .S(net868),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_095_  (.A0(\i_ibex/cs_registers_i/mtval_q [2]),
    .A1(\i_ibex/cs_registers_i/mtval_d [2]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_096_  (.A0(\i_ibex/cs_registers_i/mtval_q [30]),
    .A1(\i_ibex/cs_registers_i/mtval_d [30]),
    .S(net868),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_097_  (.A0(\i_ibex/cs_registers_i/mtval_q [31]),
    .A1(\i_ibex/cs_registers_i/mtval_d [31]),
    .S(net866),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_098_  (.A0(\i_ibex/cs_registers_i/mtval_q [3]),
    .A1(\i_ibex/cs_registers_i/mtval_d [3]),
    .S(net866),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_099_  (.A0(\i_ibex/cs_registers_i/mtval_q [4]),
    .A1(\i_ibex/cs_registers_i/mtval_d [4]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_100_  (.A0(\i_ibex/cs_registers_i/mtval_q [5]),
    .A1(\i_ibex/cs_registers_i/mtval_d [5]),
    .S(net865),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_101_  (.A0(\i_ibex/cs_registers_i/mtval_q [6]),
    .A1(\i_ibex/cs_registers_i/mtval_d [6]),
    .S(net864),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_102_  (.A0(\i_ibex/cs_registers_i/mtval_q [7]),
    .A1(\i_ibex/cs_registers_i/mtval_d [7]),
    .S(net865),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_103_  (.A0(\i_ibex/cs_registers_i/mtval_q [8]),
    .A1(\i_ibex/cs_registers_i/mtval_d [8]),
    .S(net865),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtval_csr/_104_  (.A0(\i_ibex/cs_registers_i/mtval_q [9]),
    .A1(\i_ibex/cs_registers_i/mtval_d [9]),
    .S(net866),
    .X(\i_ibex/cs_registers_i/u_mtval_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1387__55  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net55));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_81_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_000_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_067_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_80_clk_i_regs),
    .RESET_B(net1568),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_001_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_066_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_94_clk_i_regs),
    .RESET_B(net1568),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_065_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[12]_reg  (.CLK(clknet_leaf_62_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_064_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1531),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_004_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_063_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[14]_reg  (.CLK(clknet_leaf_62_clk_i_regs),
    .RESET_B(net1570),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_062_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1531),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_006_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_061_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[16]_reg  (.CLK(clknet_leaf_34_clk_i_regs),
    .RESET_B(net1634),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_060_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[17]_reg  (.CLK(clknet_leaf_40_clk_i_regs),
    .RESET_B(net1605),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_059_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[18]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1635),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_009_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_058_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1634),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_010_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_057_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_77_clk_i_regs),
    .RESET_B(net1547),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_056_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[20]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1634),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_055_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[21]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1635),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_013_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_054_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_35_clk_i_regs),
    .RESET_B(net1633),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_014_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_053_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_35_clk_i_regs),
    .RESET_B(net1634),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_052_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[24]_reg  (.CLK(clknet_leaf_34_clk_i_regs),
    .RESET_B(net1634),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_051_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_35_clk_i_regs),
    .RESET_B(net1633),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_017_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_050_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_31_clk_i_regs),
    .RESET_B(net1633),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_049_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_41_clk_i_regs),
    .RESET_B(net1606),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_048_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[28]_reg  (.CLK(clknet_leaf_33_clk_i_regs),
    .RESET_B(net1592),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_047_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_41_clk_i_regs),
    .RESET_B(net1605),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_021_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_046_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_77_clk_i_regs),
    .RESET_B(net1538),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_045_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[30]_reg  (.CLK(clknet_leaf_37_clk_i_regs),
    .RESET_B(net1635),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_044_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_94_clk_i_regs),
    .RESET_B(net1546),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_024_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_043_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_80_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_042_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_77_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_041_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_78_clk_i_regs),
    .RESET_B(net1570),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_040_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_78_clk_i_regs),
    .RESET_B(net1545),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_039_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_81_clk_i_regs),
    .RESET_B(net1569),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_038_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_78_clk_i_regs),
    .RESET_B(net1570),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_037_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtval_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_94_clk_i_regs),
    .RESET_B(net1567),
    .D(\i_ibex/cs_registers_i/u_mtval_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtval_csr/_036_ ),
    .Q(\i_ibex/cs_registers_i/mtval_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout830 (.X(net830),
    .A(net834),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout829 (.X(net829),
    .A(net830),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_072_  (.A(\i_ibex/cs_registers_i/u_mtvec_csr/_000_ ),
    .B(net894),
    .Y(\i_ibex/cs_registers_i/u_mtvec_csr/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/cs_registers_i/u_mtvec_csr/_073_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net381),
    .A2(net893),
    .Y(\i_ibex/cs_registers_i/u_mtvec_csr/_001_ ),
    .B1(\i_ibex/cs_registers_i/u_mtvec_csr/_033_ ));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_074_  (.A0(\i_ibex/csr_mtvec [10]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [10]),
    .S(net894),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_075_  (.A0(\i_ibex/csr_mtvec [11]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [11]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_076_  (.A0(\i_ibex/csr_mtvec [12]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [12]),
    .S(net894),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_077_  (.A0(\i_ibex/csr_mtvec [13]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [13]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_078_  (.A0(\i_ibex/csr_mtvec [14]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [14]),
    .S(net894),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_079_  (.A0(\i_ibex/csr_mtvec [15]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [15]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_080_  (.A0(\i_ibex/csr_mtvec [16]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [16]),
    .S(net896),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_081_  (.A0(\i_ibex/csr_mtvec [17]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [17]),
    .S(net896),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_083_  (.A0(\i_ibex/csr_mtvec [18]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [18]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_084_  (.A0(\i_ibex/csr_mtvec [19]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [19]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_085_  (.A0(\i_ibex/csr_mtvec [1]),
    .A1(net47),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_086_  (.A0(\i_ibex/csr_mtvec [20]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [20]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_087_  (.A0(\i_ibex/csr_mtvec [21]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [21]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_088_  (.A0(\i_ibex/csr_mtvec [22]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [22]),
    .S(net896),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_089_  (.A0(\i_ibex/csr_mtvec [23]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [23]),
    .S(net896),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_090_  (.A0(\i_ibex/csr_mtvec [24]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [24]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_091_  (.A0(\i_ibex/csr_mtvec [25]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [25]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_092_  (.A0(\i_ibex/csr_mtvec [26]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [26]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout827 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0237_ ),
    .X(net827),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_094_  (.A0(\i_ibex/csr_mtvec [27]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [27]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_095_  (.A0(\i_ibex/csr_mtvec [28]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [28]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_096_  (.A0(\i_ibex/csr_mtvec [29]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [29]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_097_  (.A0(\i_ibex/csr_mtvec [2]),
    .A1(net48),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_098_  (.A0(\i_ibex/csr_mtvec [30]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [30]),
    .S(net895),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_099_  (.A0(\i_ibex/csr_mtvec [31]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [31]),
    .S(net896),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_100_  (.A0(\i_ibex/csr_mtvec [3]),
    .A1(net49),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_101_  (.A0(\i_ibex/csr_mtvec [4]),
    .A1(net50),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_102_  (.A0(\i_ibex/csr_mtvec [5]),
    .A1(net51),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_103_  (.A0(\i_ibex/csr_mtvec [6]),
    .A1(net52),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_104_  (.A0(\i_ibex/csr_mtvec [7]),
    .A1(net53),
    .S(net893),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_105_  (.A0(\i_ibex/csr_mtvec [8]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [8]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/cs_registers_i/u_mtvec_csr/_106_  (.A0(\i_ibex/csr_mtvec [9]),
    .A1(\i_ibex/cs_registers_i/mtvec_d [9]),
    .S(net897),
    .X(\i_ibex/cs_registers_i/u_mtvec_csr/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1349__54  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net54));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[0]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1539),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_001_ ),
    .Q_N(\i_ibex/csr_mtvec [0]),
    .Q(\i_ibex/cs_registers_i/u_mtvec_csr/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[10]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1531),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_002_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_068_ ),
    .Q(\i_ibex/csr_mtvec [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[11]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1606),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_003_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_067_ ),
    .Q(\i_ibex/csr_mtvec [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[12]_reg  (.RESET_B(net1532),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_004_ ),
    .Q(\i_ibex/csr_mtvec [12]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_066_ ),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[13]_reg  (.CLK(clknet_leaf_39_clk_i_regs),
    .RESET_B(net1604),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_005_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_065_ ),
    .Q(\i_ibex/csr_mtvec [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[14]_reg  (.RESET_B(net1532),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_006_ ),
    .Q(\i_ibex/csr_mtvec [14]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_064_ ),
    .CLK(clknet_5_25__leaf_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[15]_reg  (.CLK(clknet_leaf_39_clk_i_regs),
    .RESET_B(net1595),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_007_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_063_ ),
    .Q(\i_ibex/csr_mtvec [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[16]_reg  (.CLK(clknet_5_3__leaf_clk_i_regs),
    .RESET_B(net1630),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_008_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_062_ ),
    .Q(\i_ibex/csr_mtvec [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[17]_reg  (.RESET_B(net1648),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_009_ ),
    .Q(\i_ibex/csr_mtvec [17]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_061_ ),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[18]_reg  (.RESET_B(net1648),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_010_ ),
    .Q(\i_ibex/csr_mtvec [18]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_060_ ),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[19]_reg  (.CLK(clknet_leaf_25_clk_i_regs),
    .RESET_B(net1648),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_011_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_059_ ),
    .Q(\i_ibex/csr_mtvec [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[1]_reg  (.CLK(clknet_leaf_64_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_012_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_058_ ),
    .Q(\i_ibex/csr_mtvec [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[20]_reg  (.RESET_B(net1628),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_013_ ),
    .Q(\i_ibex/csr_mtvec [20]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_057_ ),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[21]_reg  (.RESET_B(net1648),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_014_ ),
    .Q(\i_ibex/csr_mtvec [21]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_056_ ),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[22]_reg  (.CLK(clknet_leaf_32_clk_i_regs),
    .RESET_B(net1630),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_015_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_055_ ),
    .Q(\i_ibex/csr_mtvec [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[23]_reg  (.CLK(clknet_leaf_25_clk_i_regs),
    .RESET_B(net1629),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_016_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_054_ ),
    .Q(\i_ibex/csr_mtvec [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[24]_reg  (.RESET_B(net1645),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_017_ ),
    .Q(\i_ibex/csr_mtvec [24]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_053_ ),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[25]_reg  (.CLK(clknet_leaf_27_clk_i_regs),
    .RESET_B(net1648),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_018_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_052_ ),
    .Q(\i_ibex/csr_mtvec [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[26]_reg  (.CLK(clknet_leaf_25_clk_i_regs),
    .RESET_B(net1648),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_019_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_051_ ),
    .Q(\i_ibex/csr_mtvec [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[27]_reg  (.CLK(clknet_leaf_39_clk_i_regs),
    .RESET_B(net1595),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_020_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_050_ ),
    .Q(\i_ibex/csr_mtvec [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[28]_reg  (.RESET_B(net1595),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_021_ ),
    .Q(\i_ibex/csr_mtvec [28]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_049_ ),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[29]_reg  (.CLK(clknet_leaf_40_clk_i_regs),
    .RESET_B(net1604),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_022_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_048_ ),
    .Q(\i_ibex/csr_mtvec [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[2]_reg  (.CLK(clknet_leaf_65_clk_i_regs),
    .RESET_B(net1536),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_023_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_047_ ),
    .Q(\i_ibex/csr_mtvec [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[30]_reg  (.RESET_B(net1628),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_024_ ),
    .Q(\i_ibex/csr_mtvec [30]),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_046_ ),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[31]_reg  (.CLK(clknet_leaf_32_clk_i_regs),
    .RESET_B(net1596),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_025_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_045_ ),
    .Q(\i_ibex/csr_mtvec [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[3]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1536),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_026_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_044_ ),
    .Q(\i_ibex/csr_mtvec [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[4]_reg  (.CLK(clknet_leaf_63_clk_i_regs),
    .RESET_B(net1537),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_027_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_043_ ),
    .Q(\i_ibex/csr_mtvec [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[5]_reg  (.CLK(clknet_leaf_60_clk_i_regs),
    .RESET_B(net1530),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_028_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_042_ ),
    .Q(\i_ibex/csr_mtvec [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[6]_reg  (.CLK(clknet_leaf_68_clk_i_regs),
    .RESET_B(net1535),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_029_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_041_ ),
    .Q(\i_ibex/csr_mtvec [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[7]_reg  (.CLK(clknet_leaf_65_clk_i_regs),
    .RESET_B(net1536),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_030_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_040_ ),
    .Q(\i_ibex/csr_mtvec [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[8]_reg  (.CLK(clknet_leaf_40_clk_i_regs),
    .RESET_B(net1604),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_031_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_039_ ),
    .Q(\i_ibex/csr_mtvec [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/cs_registers_i/u_mtvec_csr/rd_data_o[9]_reg  (.CLK(clknet_leaf_43_clk_i_regs),
    .RESET_B(net1531),
    .D(\i_ibex/cs_registers_i/u_mtvec_csr/_032_ ),
    .Q_N(\i_ibex/cs_registers_i/u_mtvec_csr/_038_ ),
    .Q(\i_ibex/csr_mtvec [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/_1_  (.A(net254),
    .B(net255),
    .Y(\i_ibex/ex_valid ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/_1__254  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net254));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(net827),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout825 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0260_ ),
    .X(net825),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout824 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0260_ ),
    .X(net824),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout823 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0355_ ),
    .X(net823),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout822 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0366_ ),
    .X(net822),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout821 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0366_ ),
    .X(net821),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout820 (.X(net820),
    .A(net821),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1356_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0597_ ),
    .A(net1291),
    .VSS(VSS));
 sg13g2_buf_8 fanout819 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_158_ ),
    .X(net819),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout818 (.X(net818),
    .A(net819),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1359_  (.A(\i_ibex/alu_operator_ex [5]),
    .B_N(\i_ibex/alu_operator_ex [4]),
    .Y(\i_ibex/ex_block_i/alu_i/_0600_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1360_  (.A(net322),
    .B(net621),
    .Y(\i_ibex/ex_block_i/alu_i/_0601_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout817 (.X(net817),
    .A(net819),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/ex_block_i/alu_i/_1362_  (.Y(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .A(net1289),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1363_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0601_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0600_ ),
    .A1(net622),
    .Y(\i_ibex/ex_block_i/alu_i/_0604_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0597_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1364_  (.Y(\i_ibex/ex_block_i/alu_i/_0605_ ),
    .B(net1291),
    .A_N(net621),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_1365_  (.B(\i_ibex/alu_operator_ex [4]),
    .C(net621),
    .Y(\i_ibex/ex_block_i/alu_i/_0606_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/alu_operator_ex [5]));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1366_  (.X(\i_ibex/ex_block_i/alu_i/_0607_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0605_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0606_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1367_  (.Y(\i_ibex/ex_block_i/alu_i/_0608_ ),
    .A(\i_ibex/alu_operator_ex [4]),
    .B(\i_ibex/alu_operator_ex [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout816 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_158_ ),
    .X(net816),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1369_  (.Y(\i_ibex/ex_block_i/alu_i/_0610_ ),
    .B(net1293),
    .A_N(net323),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/ex_block_i/alu_i/_1370_  (.A(\i_ibex/ex_block_i/alu_i/_0604_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0607_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0608_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0611_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0610_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1371_  (.Y(\i_ibex/ex_block_i/alu_i/_0612_ ),
    .B(\i_ibex/alu_operator_ex [4]),
    .A_N(\i_ibex/alu_operator_ex [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout815 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_158_ ),
    .X(net815),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1373_  (.Y(\i_ibex/ex_block_i/alu_i/_0614_ ),
    .A(net621),
    .B(net1291),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/ex_block_i/alu_i/_1374_  (.A(\i_ibex/ex_block_i/alu_i/_0612_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0610_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0614_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0615_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1375_  (.Y(\i_ibex/ex_block_i/alu_i/_0616_ ),
    .B(net1289),
    .A_N(net622),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1376_  (.Y(\i_ibex/ex_block_i/alu_i/_0617_ ),
    .B(\i_ibex/alu_operator_ex [5]),
    .A_N(net1289),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/ex_block_i/alu_i/_1377_  (.A(net324),
    .B(\i_ibex/alu_operator_ex [4]),
    .C(net1291),
    .D(net1293),
    .X(\i_ibex/ex_block_i/alu_i/_0618_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1378_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0616_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0617_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0619_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0618_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1379_  (.A2(\i_ibex/ex_block_i/alu_i/_0615_ ),
    .A1(net1288),
    .B1(\i_ibex/ex_block_i/alu_i/_0619_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0620_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1380_  (.A(\i_ibex/ex_block_i/alu_i/_0611_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0620_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0621_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout814 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_169_ ),
    .X(net814),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout813 (.X(net813),
    .A(net814),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout812 (.X(net812),
    .A(net814),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout811 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_169_ ),
    .X(net811),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1385_  (.Y(\i_ibex/ex_block_i/alu_i/_0626_ ),
    .A(net532),
    .B(\i_ibex/alu_operand_b_ex [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1386_  (.Y(\i_ibex/ex_block_i/alu_i/_0627_ ),
    .A(net596),
    .B(\i_ibex/ex_block_i/alu_i/_0626_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout810 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_169_ ),
    .X(net810),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout809 (.A(net54),
    .X(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout808 (.A(net809),
    .X(net808),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1394_  (.A(\i_ibex/alu_operand_b_ex [26]),
    .B(net603),
    .Y(\i_ibex/ex_block_i/alu_i/_0635_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1395_  (.A(net56),
    .B(\i_ibex/ex_block_i/alu_i/_0635_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0636_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1396_  (.Y(\i_ibex/ex_block_i/alu_i/_0637_ ),
    .A(net57),
    .B(\i_ibex/ex_block_i/alu_i/_0636_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1397_  (.Y(\i_ibex/ex_block_i/alu_i/_0638_ ),
    .A(net793),
    .B(\i_ibex/ex_block_i/alu_i/_0637_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1398_  (.B1(\i_ibex/ex_block_i/alu_i/_0638_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0639_ ),
    .VSS(VSS),
    .A1(net801),
    .A2(\i_ibex/ex_block_i/alu_i/_0627_ ));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1400_  (.Y(\i_ibex/ex_block_i/alu_i/_0641_ ),
    .A(net529),
    .B(\i_ibex/alu_operand_b_ex [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1401_  (.Y(\i_ibex/ex_block_i/alu_i/_0642_ ),
    .A(net596),
    .B(\i_ibex/ex_block_i/alu_i/_0641_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1402_  (.A(\i_ibex/alu_operand_b_ex [25]),
    .B(net603),
    .Y(\i_ibex/ex_block_i/alu_i/_0643_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1403_  (.A(net58),
    .B(\i_ibex/ex_block_i/alu_i/_0643_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0644_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1404_  (.Y(\i_ibex/ex_block_i/alu_i/_0645_ ),
    .A(net59),
    .B(\i_ibex/ex_block_i/alu_i/_0644_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1405_  (.Y(\i_ibex/ex_block_i/alu_i/_0646_ ),
    .A(net793),
    .B(\i_ibex/ex_block_i/alu_i/_0645_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1406_  (.B1(\i_ibex/ex_block_i/alu_i/_0646_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0647_ ),
    .VSS(VSS),
    .A1(net801),
    .A2(\i_ibex/ex_block_i/alu_i/_0642_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1407_  (.A(\i_ibex/alu_operand_b_ex [24]),
    .B(net602),
    .Y(\i_ibex/ex_block_i/alu_i/_0648_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1408_  (.A(net60),
    .B(\i_ibex/ex_block_i/alu_i/_0648_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0649_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1409_  (.Y(\i_ibex/ex_block_i/alu_i/_0650_ ),
    .A(net61),
    .B(\i_ibex/ex_block_i/alu_i/_0649_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout802 (.A(net809),
    .X(net802),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1411_  (.Y(\i_ibex/ex_block_i/alu_i/_0652_ ),
    .A(net527),
    .B(\i_ibex/alu_operand_b_ex [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1412_  (.Y(\i_ibex/ex_block_i/alu_i/_0653_ ),
    .A(net596),
    .B(\i_ibex/ex_block_i/alu_i/_0652_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1413_  (.A(net801),
    .B(\i_ibex/ex_block_i/alu_i/_0653_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0654_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1414_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0654_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0655_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0650_ ),
    .A1(net793));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1415_  (.A(\i_ibex/alu_operand_b_ex [23]),
    .B(net602),
    .Y(\i_ibex/ex_block_i/alu_i/_0656_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1416_  (.A(net62),
    .B(\i_ibex/ex_block_i/alu_i/_0656_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0657_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1417_  (.Y(\i_ibex/ex_block_i/alu_i/_0658_ ),
    .A(net63),
    .B(\i_ibex/ex_block_i/alu_i/_0657_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1419_  (.Y(\i_ibex/ex_block_i/alu_i/_0660_ ),
    .A(net593),
    .B(\i_ibex/alu_operand_b_ex [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1420_  (.Y(\i_ibex/ex_block_i/alu_i/_0661_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0660_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1421_  (.A(net800),
    .B(\i_ibex/ex_block_i/alu_i/_0661_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0662_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1422_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0662_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0663_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0658_ ),
    .A1(net806));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1423_  (.A(\i_ibex/ex_block_i/alu_i/_0655_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0663_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0664_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1424_  (.X(\i_ibex/ex_block_i/alu_i/_0665_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0639_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0647_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0664_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1426_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0667_ ),
    .A(\i_ibex/alu_operand_b_ex [20]),
    .VSS(VSS));
 sg13g2_or4_2 \i_ibex/ex_block_i/alu_i/_1427_  (.A(\i_ibex/ex_block_i/alu_i/_0604_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0607_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0608_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0610_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1428_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0619_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0669_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0615_ ),
    .A1(net1288));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1429_  (.Y(\i_ibex/ex_block_i/alu_i/_0670_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0669_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1430_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0667_ ),
    .A2(net1159),
    .Y(\i_ibex/ex_block_i/alu_i/_0671_ ),
    .B1(net64));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1431_  (.Y(\i_ibex/ex_block_i/alu_i/_0672_ ),
    .A(net65),
    .B(\i_ibex/ex_block_i/alu_i/_0671_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1433_  (.Y(\i_ibex/ex_block_i/alu_i/_0674_ ),
    .A(net578),
    .B(\i_ibex/alu_operand_b_ex [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1434_  (.Y(\i_ibex/ex_block_i/alu_i/_0675_ ),
    .A(net595),
    .B(\i_ibex/ex_block_i/alu_i/_0674_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1435_  (.A(net800),
    .B(\i_ibex/ex_block_i/alu_i/_0675_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0676_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1436_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0676_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0677_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0672_ ),
    .A1(net807));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(net809),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout797 (.A(net55),
    .X(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1439_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0680_ ),
    .A(\i_ibex/alu_operand_b_ex [22]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1440_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0680_ ),
    .A2(net1159),
    .Y(\i_ibex/ex_block_i/alu_i/_0681_ ),
    .B1(net66));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1441_  (.Y(\i_ibex/ex_block_i/alu_i/_0682_ ),
    .A(net67),
    .B(\i_ibex/ex_block_i/alu_i/_0681_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1443_  (.Y(\i_ibex/ex_block_i/alu_i/_0684_ ),
    .A(net591),
    .B(\i_ibex/alu_operand_b_ex [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1444_  (.Y(\i_ibex/ex_block_i/alu_i/_0685_ ),
    .A(net599),
    .B(\i_ibex/ex_block_i/alu_i/_0684_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/ex_block_i/alu_i/_1445_  (.A(net802),
    .B(\i_ibex/ex_block_i/alu_i/_0685_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0686_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1446_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0686_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0687_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0682_ ),
    .A1(net794));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1447_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0688_ ),
    .A(\i_ibex/alu_operand_b_ex [21]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1448_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0688_ ),
    .A2(net1159),
    .Y(\i_ibex/ex_block_i/alu_i/_0689_ ),
    .B1(net68));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1449_  (.Y(\i_ibex/ex_block_i/alu_i/_0690_ ),
    .A(net69),
    .B(\i_ibex/ex_block_i/alu_i/_0689_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1451_  (.Y(\i_ibex/ex_block_i/alu_i/_0692_ ),
    .A(net580),
    .B(\i_ibex/alu_operand_b_ex [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1452_  (.Y(\i_ibex/ex_block_i/alu_i/_0693_ ),
    .A(net595),
    .B(\i_ibex/ex_block_i/alu_i/_0692_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1453_  (.A(net800),
    .B(\i_ibex/ex_block_i/alu_i/_0693_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0694_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1454_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0694_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0690_ ),
    .A1(net794));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1456_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0697_ ),
    .A(\i_ibex/alu_operand_b_ex [19]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1457_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0697_ ),
    .A2(net1159),
    .Y(\i_ibex/ex_block_i/alu_i/_0698_ ),
    .B1(net70));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1458_  (.Y(\i_ibex/ex_block_i/alu_i/_0699_ ),
    .A(net71),
    .B(\i_ibex/ex_block_i/alu_i/_0698_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1460_  (.Y(\i_ibex/ex_block_i/alu_i/_0701_ ),
    .A(net576),
    .B(\i_ibex/alu_operand_b_ex [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1461_  (.Y(\i_ibex/ex_block_i/alu_i/_0702_ ),
    .A(net595),
    .B(\i_ibex/ex_block_i/alu_i/_0701_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1462_  (.A(net801),
    .B(\i_ibex/ex_block_i/alu_i/_0702_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0703_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1463_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0703_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0704_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0699_ ),
    .A1(net794));
 sg13g2_or4_1 \i_ibex/ex_block_i/alu_i/_1464_  (.A(net452),
    .B(\i_ibex/ex_block_i/alu_i/_0687_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0704_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0705_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1465_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0706_ ),
    .A(net803),
    .VSS(VSS));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout789 (.X(net789),
    .A(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1470_  (.Y(\i_ibex/ex_block_i/alu_i/_0711_ ),
    .A(net551),
    .B(\i_ibex/alu_operand_b_ex [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1471_  (.Y(\i_ibex/ex_block_i/alu_i/_0712_ ),
    .A(net1156),
    .B(\i_ibex/ex_block_i/alu_i/_0711_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1472_  (.Y(\i_ibex/ex_block_i/alu_i/_0713_ ),
    .A(net1495),
    .B(\i_ibex/ex_block_i/alu_i/_0712_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1473_  (.A(\i_ibex/alu_operand_b_ex [7]),
    .B(net603),
    .Y(\i_ibex/ex_block_i/alu_i/_0714_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1474_  (.A(net72),
    .B(\i_ibex/ex_block_i/alu_i/_0714_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0715_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1475_  (.Y(\i_ibex/ex_block_i/alu_i/_0716_ ),
    .A(net73),
    .B(\i_ibex/ex_block_i/alu_i/_0715_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1476_  (.Y(\i_ibex/ex_block_i/alu_i/_0717_ ),
    .A(net805),
    .B(\i_ibex/ex_block_i/alu_i/_0716_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1477_  (.A(net74),
    .B(net75),
    .X(\i_ibex/ex_block_i/alu_i/_0718_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1479_  (.A(net547),
    .B(\i_ibex/alu_operand_b_ex [5]),
    .X(\i_ibex/ex_block_i/alu_i/_0720_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/ex_block_i/alu_i/_1480_  (.A(net76),
    .B(\i_ibex/ex_block_i/alu_i/_0611_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0620_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0721_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(net797),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(\i_ibex/priv_mode_id [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1483_  (.A(net795),
    .B_N(net546),
    .Y(\i_ibex/ex_block_i/alu_i/_0724_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1484_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net804),
    .A2(net77),
    .Y(\i_ibex/ex_block_i/alu_i/_0725_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0724_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1485_  (.A(\i_ibex/alu_operand_b_ex [5]),
    .B(net596),
    .C(\i_ibex/ex_block_i/alu_i/_0725_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0726_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1486_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1152),
    .C1(\i_ibex/ex_block_i/alu_i/_0726_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0720_ ),
    .A1(net805),
    .Y(\i_ibex/ex_block_i/alu_i/_0727_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0718_ ));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(\i_ibex/priv_mode_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1488_  (.A(\i_ibex/alu_operand_b_ex [6]),
    .B(net603),
    .Y(\i_ibex/ex_block_i/alu_i/_0729_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(\i_ibex/debug_mode ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1490_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/alu_operand_b_ex [6]),
    .A2(net602),
    .Y(\i_ibex/ex_block_i/alu_i/_0731_ ),
    .B1(net549));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1491_  (.A(net800),
    .B(\i_ibex/ex_block_i/alu_i/_0731_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0732_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1492_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0733_ ),
    .A(net78),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1493_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0734_ ),
    .A(net79),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1494_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0733_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0734_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0735_ ),
    .B1(net1495));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1495_  (.A(\i_ibex/ex_block_i/alu_i/_0729_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0732_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0735_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0736_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1496_  (.A(\i_ibex/ex_block_i/alu_i/_0727_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0736_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0737_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1497_  (.A0(net549),
    .A1(net80),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_0738_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(\i_ibex/instr_is_compressed_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1499_  (.B(net81),
    .C(net82),
    .A(net796),
    .Y(\i_ibex/ex_block_i/alu_i/_0740_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1500_  (.B(\i_ibex/alu_operand_b_ex [6]),
    .C(net1152),
    .A(net549),
    .Y(\i_ibex/ex_block_i/alu_i/_0741_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1501_  (.Y(\i_ibex/ex_block_i/alu_i/_0742_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0740_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0741_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1502_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0738_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0729_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0743_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0742_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1503_  (.A(\i_ibex/ex_block_i/alu_i/_0737_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_0743_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0744_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1504_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0745_ ),
    .A(\i_ibex/alu_operand_b_ex [5]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1505_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0745_ ),
    .A2(net1157),
    .Y(\i_ibex/ex_block_i/alu_i/_0746_ ),
    .B1(net83));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1506_  (.Y(\i_ibex/ex_block_i/alu_i/_0747_ ),
    .A(net84),
    .B(\i_ibex/ex_block_i/alu_i/_0746_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1507_  (.Y(\i_ibex/ex_block_i/alu_i/_0748_ ),
    .A(net546),
    .B(\i_ibex/alu_operand_b_ex [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1508_  (.Y(\i_ibex/ex_block_i/alu_i/_0749_ ),
    .A(net597),
    .B(\i_ibex/ex_block_i/alu_i/_0748_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1509_  (.A(net796),
    .B(\i_ibex/ex_block_i/alu_i/_0749_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0750_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1510_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net792),
    .A2(\i_ibex/ex_block_i/alu_i/_0747_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0751_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0750_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1511_  (.B1(\i_ibex/ex_block_i/alu_i/_0734_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0752_ ),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_b_ex [6]),
    .A2(net599));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1512_  (.Y(\i_ibex/ex_block_i/alu_i/_0753_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0733_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0752_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1513_  (.Y(\i_ibex/ex_block_i/alu_i/_0754_ ),
    .A(net548),
    .B(\i_ibex/alu_operand_b_ex [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1514_  (.Y(\i_ibex/ex_block_i/alu_i/_0755_ ),
    .A(net597),
    .B(\i_ibex/ex_block_i/alu_i/_0754_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1515_  (.A(net794),
    .B(\i_ibex/ex_block_i/alu_i/_0755_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0756_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1516_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0756_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0757_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0753_ ),
    .A1(net800));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1517_  (.A(\i_ibex/ex_block_i/alu_i/_0751_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0757_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0758_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout782 (.A(net783),
    .X(net782),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1519_  (.A0(net542),
    .A1(net85),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_0760_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(net783),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1521_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0669_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0762_ ),
    .B1(\i_ibex/alu_operand_b_ex [3]));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1522_  (.Y(\i_ibex/ex_block_i/alu_i/_0763_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0760_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0762_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1523_  (.B(net86),
    .C(net87),
    .A(net790),
    .Y(\i_ibex/ex_block_i/alu_i/_0764_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1524_  (.A(net542),
    .B(\i_ibex/alu_operand_b_ex [3]),
    .X(\i_ibex/ex_block_i/alu_i/_0765_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1525_  (.Y(\i_ibex/ex_block_i/alu_i/_0766_ ),
    .A(net1153),
    .B(\i_ibex/ex_block_i/alu_i/_0765_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1526_  (.X(\i_ibex/ex_block_i/alu_i/_0767_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0763_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0764_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0766_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1527_  (.A(net88),
    .B(net89),
    .X(\i_ibex/ex_block_i/alu_i/_0768_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout780 (.A(\i_ibex/id_stage_i/imm_u_type [12]),
    .X(net780),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1530_  (.A(net545),
    .B(\i_ibex/alu_operand_b_ex [4]),
    .X(\i_ibex/ex_block_i/alu_i/_0771_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1531_  (.A(net790),
    .B_N(net544),
    .Y(\i_ibex/ex_block_i/alu_i/_0772_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1532_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net795),
    .A2(net90),
    .Y(\i_ibex/ex_block_i/alu_i/_0773_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0772_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1533_  (.A(\i_ibex/alu_operand_b_ex [4]),
    .B(net596),
    .C(\i_ibex/ex_block_i/alu_i/_0773_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0774_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1534_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1152),
    .C1(\i_ibex/ex_block_i/alu_i/_0774_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0771_ ),
    .A1(net796),
    .Y(\i_ibex/ex_block_i/alu_i/_0775_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0768_ ));
 sg13g2_buf_2 fanout778 (.A(net780),
    .X(net778),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1536_  (.A0(net540),
    .A1(net91),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_0777_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout777 (.A(\i_ibex/id_stage_i/imm_u_type [13]),
    .X(net777),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1538_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0669_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0779_ ),
    .B1(\i_ibex/alu_operand_b_ex [2]));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1539_  (.A(net540),
    .B(\i_ibex/alu_operand_b_ex [2]),
    .X(\i_ibex/ex_block_i/alu_i/_0780_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1540_  (.X(\i_ibex/ex_block_i/alu_i/_0781_ ),
    .A(net801),
    .B(net92),
    .C(net93),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1541_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1153),
    .C1(\i_ibex/ex_block_i/alu_i/_0781_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0780_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0777_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0782_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0779_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1542_  (.Y(\i_ibex/ex_block_i/alu_i/_0783_ ),
    .A(net540),
    .B(\i_ibex/alu_operand_b_ex [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1543_  (.Y(\i_ibex/ex_block_i/alu_i/_0784_ ),
    .A(net1157),
    .B(\i_ibex/ex_block_i/alu_i/_0783_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1544_  (.Y(\i_ibex/ex_block_i/alu_i/_0785_ ),
    .A(net1496),
    .B(\i_ibex/ex_block_i/alu_i/_0784_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_1545_  (.A(net94),
    .B(net95),
    .C(\i_ibex/ex_block_i/alu_i/_0779_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0786_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1546_  (.B1(net96),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0787_ ),
    .VSS(VSS),
    .A1(net97),
    .A2(\i_ibex/ex_block_i/alu_i/_0779_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1547_  (.B(\i_ibex/ex_block_i/alu_i/_0786_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0787_ ),
    .A(net804),
    .Y(\i_ibex/ex_block_i/alu_i/_0788_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1549_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0790_ ),
    .A(net526),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1550_  (.A(net98),
    .B(net99),
    .Y(\i_ibex/ex_block_i/alu_i/_0791_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout775 (.A(net777),
    .X(net775),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1552_  (.A(net799),
    .B(net536),
    .Y(\i_ibex/ex_block_i/alu_i/_0793_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1553_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net790),
    .A2(\i_ibex/ex_block_i/alu_i/_0791_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0794_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0793_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1554_  (.A(\i_ibex/ex_block_i/alu_i/_0790_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0794_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0795_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout774 (.A(net777),
    .X(net774),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout773 (.A(\i_ibex/id_stage_i/imm_u_type [14]),
    .X(net773),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1557_  (.Y(\i_ibex/ex_block_i/alu_i/_0798_ ),
    .B(net488),
    .A_N(net101),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1558_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net100),
    .A2(\i_ibex/ex_block_i/alu_i/_0798_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0799_ ),
    .B1(net102));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1559_  (.A(net100),
    .B(\i_ibex/ex_block_i/alu_i/_0798_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0800_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1560_  (.B1(net790),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0801_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0799_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0800_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1561_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0802_ ),
    .A(net488),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_1562_  (.A(net803),
    .B(net535),
    .C(net1052),
    .X(\i_ibex/ex_block_i/alu_i/_0803_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1563_  (.A(net535),
    .B(net488),
    .X(\i_ibex/ex_block_i/alu_i/_0804_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1564_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0805_ ),
    .A(net103),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1565_  (.B(net104),
    .C(net105),
    .A(net100),
    .Y(\i_ibex/ex_block_i/alu_i/_0806_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1566_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net100),
    .A2(net106),
    .Y(\i_ibex/ex_block_i/alu_i/_0807_ ),
    .B1(net107));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1567_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0805_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0806_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0808_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0807_ ));
 sg13g2_mux2_2 \i_ibex/ex_block_i/alu_i/_1568_  (.A0(\i_ibex/ex_block_i/alu_i/_0804_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0808_ ),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_0809_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1569_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0801_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0803_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0810_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0809_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1570_  (.B1(net108),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0811_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0790_ ),
    .A2(net109));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1571_  (.Y(\i_ibex/ex_block_i/alu_i/_0812_ ),
    .A(net536),
    .B(\i_ibex/ex_block_i/alu_i/_0790_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1572_  (.A0(\i_ibex/ex_block_i/alu_i/_0811_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0812_ ),
    .S(net1495),
    .X(\i_ibex/ex_block_i/alu_i/_0813_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1573_  (.B1(\i_ibex/ex_block_i/alu_i/_0813_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0814_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0795_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0810_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1574_  (.Y(\i_ibex/ex_block_i/alu_i/_0815_ ),
    .A(\i_ibex/alu_operand_b_ex [1]),
    .B(\i_ibex/ex_block_i/alu_i/_0804_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_1575_  (.Y(\i_ibex/ex_block_i/alu_i/_0816_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0815_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_0793_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0791_ ),
    .A1(net789),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1576_  (.Y(\i_ibex/ex_block_i/alu_i/_0817_ ),
    .A(net536),
    .B(net526),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1577_  (.B(net110),
    .C(net111),
    .A(net789),
    .Y(\i_ibex/ex_block_i/alu_i/_0818_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1578_  (.B1(\i_ibex/ex_block_i/alu_i/_0818_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0819_ ),
    .VSS(VSS),
    .A1(net787),
    .A2(\i_ibex/ex_block_i/alu_i/_0817_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1579_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0809_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0816_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0820_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0819_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1580_  (.Y(\i_ibex/ex_block_i/alu_i/_0821_ ),
    .A(net602),
    .B(\i_ibex/ex_block_i/alu_i/_0820_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1581_  (.B1(\i_ibex/ex_block_i/alu_i/_0821_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0822_ ),
    .VSS(VSS),
    .A1(net597),
    .A2(\i_ibex/ex_block_i/alu_i/_0814_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1582_  (.A2(\i_ibex/ex_block_i/alu_i/_0788_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0785_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0822_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0823_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_1583_  (.B(\i_ibex/ex_block_i/alu_i/_0775_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0782_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0767_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0824_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0823_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1584_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0825_ ),
    .A(\i_ibex/alu_operand_b_ex [4]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1585_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0825_ ),
    .A2(net1157),
    .Y(\i_ibex/ex_block_i/alu_i/_0826_ ),
    .B1(net112));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1586_  (.Y(\i_ibex/ex_block_i/alu_i/_0827_ ),
    .A(net113),
    .B(\i_ibex/ex_block_i/alu_i/_0826_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1587_  (.Y(\i_ibex/ex_block_i/alu_i/_0828_ ),
    .A(net544),
    .B(\i_ibex/alu_operand_b_ex [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1588_  (.Y(\i_ibex/ex_block_i/alu_i/_0829_ ),
    .A(net595),
    .B(\i_ibex/ex_block_i/alu_i/_0828_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1589_  (.A(net801),
    .B(\i_ibex/ex_block_i/alu_i/_0829_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0830_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1590_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0830_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0831_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0827_ ),
    .A1(net794));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1591_  (.B(\i_ibex/ex_block_i/alu_i/_0764_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0766_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0763_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0832_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1592_  (.Y(\i_ibex/ex_block_i/alu_i/_0833_ ),
    .A(net542),
    .B(\i_ibex/alu_operand_b_ex [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1593_  (.Y(\i_ibex/ex_block_i/alu_i/_0834_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0833_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1594_  (.A(net793),
    .B(\i_ibex/ex_block_i/alu_i/_0834_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0835_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_1595_  (.A(net114),
    .B(net115),
    .C(\i_ibex/ex_block_i/alu_i/_0762_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0836_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1596_  (.B1(net116),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0837_ ),
    .VSS(VSS),
    .A1(net117),
    .A2(\i_ibex/ex_block_i/alu_i/_0762_ ));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1597_  (.X(\i_ibex/ex_block_i/alu_i/_0838_ ),
    .A(net801),
    .B(\i_ibex/ex_block_i/alu_i/_0836_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0837_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1598_  (.A(\i_ibex/ex_block_i/alu_i/_0832_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0835_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0838_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0839_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1599_  (.B1(\i_ibex/ex_block_i/alu_i/_0775_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0840_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0831_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0839_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1600_  (.B(\i_ibex/ex_block_i/alu_i/_0824_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0840_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0758_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0841_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1601_  (.A(\i_ibex/alu_operand_b_ex [8]),
    .B(net603),
    .Y(\i_ibex/ex_block_i/alu_i/_0842_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1602_  (.A(net118),
    .B(\i_ibex/ex_block_i/alu_i/_0842_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0843_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1603_  (.Y(\i_ibex/ex_block_i/alu_i/_0844_ ),
    .A(net119),
    .B(\i_ibex/ex_block_i/alu_i/_0843_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout772 (.A(net773),
    .X(net772),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1605_  (.Y(\i_ibex/ex_block_i/alu_i/_0846_ ),
    .A(net553),
    .B(\i_ibex/alu_operand_b_ex [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1606_  (.Y(\i_ibex/ex_block_i/alu_i/_0847_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0846_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1607_  (.A(net792),
    .B(\i_ibex/ex_block_i/alu_i/_0847_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0848_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1608_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0848_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0849_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0844_ ),
    .A1(net805));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1609_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0850_ ),
    .A(\i_ibex/alu_operand_b_ex [10]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1610_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0850_ ),
    .A2(net1156),
    .Y(\i_ibex/ex_block_i/alu_i/_0851_ ),
    .B1(net120));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1611_  (.Y(\i_ibex/ex_block_i/alu_i/_0852_ ),
    .A(net121),
    .B(\i_ibex/ex_block_i/alu_i/_0851_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout771 (.A(net773),
    .X(net771),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1613_  (.Y(\i_ibex/ex_block_i/alu_i/_0854_ ),
    .A(net557),
    .B(\i_ibex/alu_operand_b_ex [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1614_  (.Y(\i_ibex/ex_block_i/alu_i/_0855_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0854_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1615_  (.A(net791),
    .B(\i_ibex/ex_block_i/alu_i/_0855_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0856_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1616_  (.A2(\i_ibex/ex_block_i/alu_i/_0852_ ),
    .A1(net805),
    .B1(\i_ibex/ex_block_i/alu_i/_0856_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0857_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout770 (.A(net773),
    .X(net770),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1618_  (.Y(\i_ibex/ex_block_i/alu_i/_0859_ ),
    .A(net554),
    .B(\i_ibex/alu_operand_b_ex [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1619_  (.Y(\i_ibex/ex_block_i/alu_i/_0860_ ),
    .A(net1156),
    .B(\i_ibex/ex_block_i/alu_i/_0859_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1620_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0861_ ),
    .A(\i_ibex/alu_operand_b_ex [9]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1621_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0861_ ),
    .A2(net1156),
    .Y(\i_ibex/ex_block_i/alu_i/_0862_ ),
    .B1(net122));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1622_  (.Y(\i_ibex/ex_block_i/alu_i/_0863_ ),
    .A(net123),
    .B(\i_ibex/ex_block_i/alu_i/_0862_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/ex_block_i/alu_i/_1623_  (.A0(\i_ibex/ex_block_i/alu_i/_0860_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0863_ ),
    .S(net788),
    .X(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1624_  (.A(\i_ibex/ex_block_i/alu_i/_0857_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0865_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1625_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0866_ ),
    .A(\i_ibex/alu_operand_b_ex [14]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1626_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0866_ ),
    .A2(net1156),
    .Y(\i_ibex/ex_block_i/alu_i/_0867_ ),
    .B1(net124));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1627_  (.Y(\i_ibex/ex_block_i/alu_i/_0868_ ),
    .A(net125),
    .B(\i_ibex/ex_block_i/alu_i/_0867_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 max_cap769 (.X(net769),
    .A(\i_ibex/id_stage_i/zimm_rs1_type [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1629_  (.Y(\i_ibex/ex_block_i/alu_i/_0870_ ),
    .A(net567),
    .B(\i_ibex/alu_operand_b_ex [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1630_  (.Y(\i_ibex/ex_block_i/alu_i/_0871_ ),
    .A(net597),
    .B(\i_ibex/ex_block_i/alu_i/_0870_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1631_  (.A(net793),
    .B(\i_ibex/ex_block_i/alu_i/_0871_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0872_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1632_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0872_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0873_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0868_ ),
    .A1(net800));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1633_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0874_ ),
    .A(\i_ibex/alu_operand_b_ex [11]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1634_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0874_ ),
    .A2(net1156),
    .Y(\i_ibex/ex_block_i/alu_i/_0875_ ),
    .B1(net126));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1635_  (.Y(\i_ibex/ex_block_i/alu_i/_0876_ ),
    .A(net127),
    .B(\i_ibex/ex_block_i/alu_i/_0875_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 max_cap768 (.A(\i_ibex/id_stage_i/zimm_rs1_type [0]),
    .X(net768),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1637_  (.Y(\i_ibex/ex_block_i/alu_i/_0878_ ),
    .A(net558),
    .B(\i_ibex/alu_operand_b_ex [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1638_  (.Y(\i_ibex/ex_block_i/alu_i/_0879_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0878_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1639_  (.A(net791),
    .B(\i_ibex/ex_block_i/alu_i/_0879_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0880_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1640_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0880_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0881_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0876_ ),
    .A1(net796));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1641_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0882_ ),
    .A(\i_ibex/alu_operand_b_ex [13]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1642_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0882_ ),
    .A2(net1156),
    .Y(\i_ibex/ex_block_i/alu_i/_0883_ ),
    .B1(net128));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1643_  (.Y(\i_ibex/ex_block_i/alu_i/_0884_ ),
    .A(net129),
    .B(\i_ibex/ex_block_i/alu_i/_0883_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 max_cap767 (.X(net767),
    .A(\i_ibex/id_stage_i/zimm_rs1_type [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1645_  (.Y(\i_ibex/ex_block_i/alu_i/_0886_ ),
    .A(net565),
    .B(\i_ibex/alu_operand_b_ex [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1646_  (.Y(\i_ibex/ex_block_i/alu_i/_0887_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0886_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1647_  (.A(net791),
    .B(\i_ibex/ex_block_i/alu_i/_0887_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0888_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1648_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0888_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0884_ ),
    .A1(net795));
 sg13g2_buf_8 max_cap766 (.A(\i_ibex/id_stage_i/zimm_rs1_type [1]),
    .X(net766),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1650_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0891_ ),
    .A(net130),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1651_  (.B1(\i_ibex/ex_block_i/alu_i/_0891_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0892_ ),
    .VSS(VSS),
    .A1(net1107),
    .A2(net595));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_1652_  (.B(\i_ibex/ex_block_i/alu_i/_0892_ ),
    .A(net131),
    .X(\i_ibex/ex_block_i/alu_i/_0893_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 max_cap765 (.X(net765),
    .A(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1654_  (.Y(\i_ibex/ex_block_i/alu_i/_0895_ ),
    .A(net563),
    .B(net1107),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1655_  (.Y(\i_ibex/ex_block_i/alu_i/_0896_ ),
    .A(net598),
    .B(\i_ibex/ex_block_i/alu_i/_0895_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1656_  (.A(net791),
    .B(\i_ibex/ex_block_i/alu_i/_0896_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0897_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1657_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0897_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0898_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0893_ ),
    .A1(net795));
 sg13g2_nor4_2 \i_ibex/ex_block_i/alu_i/_1658_  (.A(\i_ibex/ex_block_i/alu_i/_0873_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0881_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0899_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0898_ ));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_1659_  (.B(\i_ibex/ex_block_i/alu_i/_0865_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0899_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0900_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/ex_block_i/alu_i/_0849_ ));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1660_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0841_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0900_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0744_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0713_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0901_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0717_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1661_  (.A0(net567),
    .A1(net132),
    .S(net799),
    .X(\i_ibex/ex_block_i/alu_i/_0902_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1662_  (.B(net1158),
    .C(\i_ibex/ex_block_i/alu_i/_0902_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0866_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0903_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1663_  (.A(\i_ibex/alu_operand_b_ex [13]),
    .B(net601),
    .Y(\i_ibex/ex_block_i/alu_i/_0904_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1664_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/alu_operand_b_ex [13]),
    .C1(\i_ibex/ex_block_i/alu_i/_0904_ ),
    .B1(net1152),
    .A1(net795),
    .Y(\i_ibex/ex_block_i/alu_i/_0905_ ),
    .A2(net133));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1665_  (.A0(net565),
    .A1(net134),
    .S(net799),
    .X(\i_ibex/ex_block_i/alu_i/_0906_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1666_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0907_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0906_ ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1667_  (.Y(\i_ibex/ex_block_i/alu_i/_0908_ ),
    .A(net558),
    .B(\i_ibex/alu_operand_b_ex [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1668_  (.B(net135),
    .C(net136),
    .A(net803),
    .Y(\i_ibex/ex_block_i/alu_i/_0909_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1669_  (.B1(\i_ibex/ex_block_i/alu_i/_0909_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0910_ ),
    .VSS(VSS),
    .A1(net799),
    .A2(\i_ibex/ex_block_i/alu_i/_0908_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1670_  (.B1(net137),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0911_ ),
    .VSS(VSS),
    .A1(net138),
    .A2(\i_ibex/ex_block_i/alu_i/_0910_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1671_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0912_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0911_ ),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1672_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net139),
    .A2(\i_ibex/ex_block_i/alu_i/_0910_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0913_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0912_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1673_  (.B(net1107),
    .C(\i_ibex/alu_operand_b_ex [11]),
    .A(net558),
    .Y(\i_ibex/ex_block_i/alu_i/_0914_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1674_  (.Y(\i_ibex/ex_block_i/alu_i/_0915_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0914_ ),
    .A_N(net562),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1675_  (.Y(\i_ibex/ex_block_i/alu_i/_0916_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0908_ ),
    .A_N(net1107),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1676_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0915_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0916_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0917_ ),
    .B1(net800));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1677_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net807),
    .A2(\i_ibex/ex_block_i/alu_i/_0913_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0918_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0917_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1678_  (.Y(\i_ibex/ex_block_i/alu_i/_0919_ ),
    .A(net558),
    .B(\i_ibex/ex_block_i/alu_i/_0874_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1679_  (.Y(\i_ibex/ex_block_i/alu_i/_0920_ ),
    .B(\i_ibex/alu_operand_b_ex [11]),
    .A_N(net140),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1680_  (.B(net141),
    .C(\i_ibex/ex_block_i/alu_i/_0920_ ),
    .A(net803),
    .Y(\i_ibex/ex_block_i/alu_i/_0921_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1681_  (.B1(\i_ibex/ex_block_i/alu_i/_0921_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0922_ ),
    .VSS(VSS),
    .A1(net799),
    .A2(\i_ibex/ex_block_i/alu_i/_0919_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1682_  (.Y(\i_ibex/ex_block_i/alu_i/_0923_ ),
    .A(net1107),
    .B(\i_ibex/ex_block_i/alu_i/_0891_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1683_  (.Y(\i_ibex/ex_block_i/alu_i/_0924_ ),
    .B(net803),
    .A_N(net142),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1684_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0922_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0923_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0925_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0924_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1685_  (.A(net1107),
    .B_N(net562),
    .Y(\i_ibex/ex_block_i/alu_i/_0926_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1686_  (.Y(\i_ibex/ex_block_i/alu_i/_0927_ ),
    .B(net1107),
    .A_N(net562),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1687_  (.B1(\i_ibex/ex_block_i/alu_i/_0927_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0928_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0926_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0922_ ));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1688_  (.A(net1495),
    .B(\i_ibex/ex_block_i/alu_i/_0928_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0929_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1689_  (.A(\i_ibex/ex_block_i/alu_i/_0922_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0923_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0930_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/ex_block_i/alu_i/_1690_  (.A(net596),
    .B(\i_ibex/ex_block_i/alu_i/_0925_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0929_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0930_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0931_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1691_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0931_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0932_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0918_ ),
    .A1(net603));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1692_  (.A2(\i_ibex/ex_block_i/alu_i/_0907_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0905_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0932_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0933_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1693_  (.Y(\i_ibex/ex_block_i/alu_i/_0934_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0906_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_0905_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1694_  (.A2(\i_ibex/ex_block_i/alu_i/_0934_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0933_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0873_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0935_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1695_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net792),
    .A2(\i_ibex/ex_block_i/alu_i/_0852_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0936_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0856_ ));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1696_  (.A(net143),
    .B(net144),
    .X(\i_ibex/ex_block_i/alu_i/_0937_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1697_  (.A(net554),
    .B(\i_ibex/alu_operand_b_ex [9]),
    .X(\i_ibex/ex_block_i/alu_i/_0938_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 max_cap764 (.X(net764),
    .A(net762),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1699_  (.A(net794),
    .B_N(net554),
    .Y(\i_ibex/ex_block_i/alu_i/_0940_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1700_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net806),
    .A2(net145),
    .Y(\i_ibex/ex_block_i/alu_i/_0941_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0940_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1701_  (.A(\i_ibex/alu_operand_b_ex [9]),
    .B(net598),
    .C(\i_ibex/ex_block_i/alu_i/_0941_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0942_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1702_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1152),
    .C1(\i_ibex/ex_block_i/alu_i/_0942_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0938_ ),
    .A1(net805),
    .Y(\i_ibex/ex_block_i/alu_i/_0943_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0937_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1703_  (.A0(net556),
    .A1(net146),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_0944_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_1704_  (.B(net1156),
    .C(\i_ibex/ex_block_i/alu_i/_0944_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0945_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/alu_operand_b_ex [10]));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1705_  (.B(net147),
    .C(net148),
    .A(net795),
    .Y(\i_ibex/ex_block_i/alu_i/_0946_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1706_  (.A(net556),
    .B(\i_ibex/alu_operand_b_ex [10]),
    .X(\i_ibex/ex_block_i/alu_i/_0947_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1707_  (.Y(\i_ibex/ex_block_i/alu_i/_0948_ ),
    .A(net1152),
    .B(\i_ibex/ex_block_i/alu_i/_0947_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1708_  (.X(\i_ibex/ex_block_i/alu_i/_0949_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0945_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0946_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0948_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1709_  (.B1(\i_ibex/ex_block_i/alu_i/_0949_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0950_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0936_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0943_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1710_  (.A0(net550),
    .A1(net149),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_0951_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1711_  (.A(net550),
    .B(\i_ibex/alu_operand_b_ex [7]),
    .X(\i_ibex/ex_block_i/alu_i/_0952_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1712_  (.X(\i_ibex/ex_block_i/alu_i/_0953_ ),
    .A(net789),
    .B(net150),
    .C(net151),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1713_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1152),
    .C1(\i_ibex/ex_block_i/alu_i/_0953_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0952_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0714_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0954_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0951_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1714_  (.A0(net553),
    .A1(net152),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_0955_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1715_  (.A(net552),
    .B(\i_ibex/alu_operand_b_ex [8]),
    .X(\i_ibex/ex_block_i/alu_i/_0956_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1716_  (.X(\i_ibex/ex_block_i/alu_i/_0957_ ),
    .A(net789),
    .B(net153),
    .C(net154),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1717_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1152),
    .C1(\i_ibex/ex_block_i/alu_i/_0957_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0956_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0842_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0958_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0955_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1718_  (.A2(net601),
    .A1(\i_ibex/alu_operand_b_ex [8]),
    .B1(net552),
    .X(\i_ibex/ex_block_i/alu_i/_0959_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1719_  (.B1(net794),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0960_ ),
    .VSS(VSS),
    .A1(net155),
    .A2(net156));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1720_  (.B1(\i_ibex/ex_block_i/alu_i/_0960_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0961_ ),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_b_ex [8]),
    .A2(net597));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1721_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1495),
    .A2(\i_ibex/ex_block_i/alu_i/_0959_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0962_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0961_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1722_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0954_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0958_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0963_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0962_ ));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1723_  (.X(\i_ibex/ex_block_i/alu_i/_0964_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0857_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0963_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1724_  (.B1(net1516),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0965_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0950_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0964_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1725_  (.B(net157),
    .C(net158),
    .A(net805),
    .Y(\i_ibex/ex_block_i/alu_i/_0966_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1726_  (.B(\i_ibex/alu_operand_b_ex [14]),
    .C(net1153),
    .A(net567),
    .Y(\i_ibex/ex_block_i/alu_i/_0967_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1727_  (.A(\i_ibex/ex_block_i/alu_i/_0966_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0967_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0968_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_1728_  (.B(\i_ibex/ex_block_i/alu_i/_0935_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0965_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0903_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0969_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0968_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1729_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0669_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0970_ ),
    .B1(\i_ibex/alu_operand_b_ex [18]));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1730_  (.A(net159),
    .B(\i_ibex/ex_block_i/alu_i/_0970_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0971_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_1731_  (.B(\i_ibex/ex_block_i/alu_i/_0971_ ),
    .A(net160),
    .X(\i_ibex/ex_block_i/alu_i/_0972_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 max_cap763 (.A(net762),
    .X(net763),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1733_  (.Y(\i_ibex/ex_block_i/alu_i/_0974_ ),
    .A(net574),
    .B(\i_ibex/alu_operand_b_ex [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1734_  (.Y(\i_ibex/ex_block_i/alu_i/_0975_ ),
    .A(net1159),
    .B(\i_ibex/ex_block_i/alu_i/_0974_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1735_  (.Y(\i_ibex/ex_block_i/alu_i/_0976_ ),
    .A(net1496),
    .B(\i_ibex/ex_block_i/alu_i/_0975_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1736_  (.B1(\i_ibex/ex_block_i/alu_i/_0976_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0977_ ),
    .VSS(VSS),
    .A1(net1496),
    .A2(\i_ibex/ex_block_i/alu_i/_0972_ ));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(\i_ibex/id_stage_i/imm_u_type [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1738_  (.Y(\i_ibex/ex_block_i/alu_i/_0979_ ),
    .A(net572),
    .B(\i_ibex/alu_operand_b_ex [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1739_  (.Y(\i_ibex/ex_block_i/alu_i/_0980_ ),
    .A(net595),
    .B(\i_ibex/ex_block_i/alu_i/_0979_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1740_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0669_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0981_ ),
    .B1(\i_ibex/alu_operand_b_ex [17]));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_1741_  (.A(net161),
    .B(net162),
    .C(\i_ibex/ex_block_i/alu_i/_0981_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0982_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1742_  (.B1(net163),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0983_ ),
    .VSS(VSS),
    .A1(net164),
    .A2(\i_ibex/ex_block_i/alu_i/_0981_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1743_  (.B(\i_ibex/ex_block_i/alu_i/_0982_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0983_ ),
    .A(net790),
    .Y(\i_ibex/ex_block_i/alu_i/_0984_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1744_  (.B1(\i_ibex/ex_block_i/alu_i/_0984_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0985_ ),
    .VSS(VSS),
    .A1(net788),
    .A2(\i_ibex/ex_block_i/alu_i/_0980_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1745_  (.Y(\i_ibex/ex_block_i/alu_i/_0986_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0977_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0985_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1746_  (.A(\i_ibex/alu_operand_b_ex [15]),
    .B(net601),
    .Y(\i_ibex/ex_block_i/alu_i/_0987_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1747_  (.A(net165),
    .B(\i_ibex/ex_block_i/alu_i/_0987_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0988_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1748_  (.Y(\i_ibex/ex_block_i/alu_i/_0989_ ),
    .A(net166),
    .B(\i_ibex/ex_block_i/alu_i/_0988_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(net763),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1750_  (.Y(\i_ibex/ex_block_i/alu_i/_0991_ ),
    .A(net569),
    .B(\i_ibex/alu_operand_b_ex [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1751_  (.Y(\i_ibex/ex_block_i/alu_i/_0992_ ),
    .A(net596),
    .B(\i_ibex/ex_block_i/alu_i/_0991_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1752_  (.A(net793),
    .B(\i_ibex/ex_block_i/alu_i/_0992_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0993_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1753_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net792),
    .A2(\i_ibex/ex_block_i/alu_i/_0989_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0994_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0993_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1754_  (.A(net789),
    .B_N(\i_ibex/alu_operand_b_ex [16]),
    .Y(\i_ibex/ex_block_i/alu_i/_0995_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1755_  (.A(\i_ibex/alu_operand_b_ex [16]),
    .B(net601),
    .Y(\i_ibex/ex_block_i/alu_i/_0996_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1756_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0995_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0996_ ),
    .B1(net595),
    .A1(net804),
    .Y(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .A2(net167));
 sg13g2_buf_16 max_cap760 (.X(net760),
    .A(net758),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1758_  (.A(net804),
    .B_N(net570),
    .Y(\i_ibex/ex_block_i/alu_i/_0999_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1759_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0999_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .A2(net168),
    .A1(net804));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1760_  (.Y(\i_ibex/ex_block_i/alu_i/_1001_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1761_  (.A(\i_ibex/ex_block_i/alu_i/_0986_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0994_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1001_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1762_  (.B1(\i_ibex/ex_block_i/alu_i/_1002_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1003_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0901_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0969_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1763_  (.B(\i_ibex/alu_operand_b_ex [18]),
    .C(net1155),
    .A(net574),
    .Y(\i_ibex/ex_block_i/alu_i/_1004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1764_  (.A0(net572),
    .A1(net169),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_1005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1765_  (.Y(\i_ibex/ex_block_i/alu_i/_1006_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1005_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0981_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1766_  (.B(net170),
    .C(net171),
    .A(net804),
    .Y(\i_ibex/ex_block_i/alu_i/_1007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1767_  (.B(\i_ibex/alu_operand_b_ex [17]),
    .C(net1155),
    .A(net571),
    .Y(\i_ibex/ex_block_i/alu_i/_1008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1768_  (.B(\i_ibex/ex_block_i/alu_i/_1007_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1008_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1006_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1769_  (.Y(\i_ibex/ex_block_i/alu_i/_1010_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0977_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1770_  (.A0(net569),
    .A1(net172),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_1011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1771_  (.A(net569),
    .B(\i_ibex/alu_operand_b_ex [15]),
    .X(\i_ibex/ex_block_i/alu_i/_1012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1772_  (.X(\i_ibex/ex_block_i/alu_i/_1013_ ),
    .A(net789),
    .B(net173),
    .C(net174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1773_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1154),
    .C1(\i_ibex/ex_block_i/alu_i/_1013_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1012_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1011_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1014_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0987_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1774_  (.B1(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1015_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1014_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1775_  (.Y(\i_ibex/ex_block_i/alu_i/_1016_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_1776_  (.B(\i_ibex/ex_block_i/alu_i/_1015_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1016_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0977_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1017_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0985_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1777_  (.A0(net573),
    .A1(net175),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_1018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1778_  (.A(net176),
    .B(net177),
    .X(\i_ibex/ex_block_i/alu_i/_1019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_1779_  (.Y(\i_ibex/ex_block_i/alu_i/_1020_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1019_ ),
    .B2(net792),
    .A2(\i_ibex/ex_block_i/alu_i/_0970_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_1780_  (.B(\i_ibex/ex_block_i/alu_i/_1010_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1017_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1004_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1021_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_1020_ ));
 sg13g2_buf_1 max_cap759 (.A(net758),
    .X(net759),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1782_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1023_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0705_ ),
    .VSS(VSS));
 sg13g2_buf_2 fanout758 (.A(\i_ibex/id_stage_i/imm_u_type [21]),
    .X(net758),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1784_  (.A(net178),
    .B(net179),
    .X(\i_ibex/ex_block_i/alu_i/_1025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1785_  (.A(net576),
    .B(\i_ibex/alu_operand_b_ex [19]),
    .X(\i_ibex/ex_block_i/alu_i/_1026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1786_  (.A(net803),
    .B_N(net575),
    .Y(\i_ibex/ex_block_i/alu_i/_1027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1787_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net790),
    .A2(net180),
    .Y(\i_ibex/ex_block_i/alu_i/_1028_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1027_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1788_  (.A(\i_ibex/alu_operand_b_ex [19]),
    .B(net597),
    .C(\i_ibex/ex_block_i/alu_i/_1028_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1789_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1154),
    .C1(\i_ibex/ex_block_i/alu_i/_1029_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1026_ ),
    .A1(net791),
    .Y(\i_ibex/ex_block_i/alu_i/_1030_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1025_ ));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1790_  (.A(net181),
    .B(net182),
    .X(\i_ibex/ex_block_i/alu_i/_1031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1791_  (.A(net577),
    .B(\i_ibex/alu_operand_b_ex [20]),
    .X(\i_ibex/ex_block_i/alu_i/_1032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1792_  (.A(net790),
    .B_N(net577),
    .Y(\i_ibex/ex_block_i/alu_i/_1033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1793_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net794),
    .A2(net183),
    .Y(\i_ibex/ex_block_i/alu_i/_1034_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1033_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1794_  (.A(\i_ibex/alu_operand_b_ex [20]),
    .B(net595),
    .C(\i_ibex/ex_block_i/alu_i/_1034_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1795_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1154),
    .C1(\i_ibex/ex_block_i/alu_i/_1035_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1032_ ),
    .A1(net793),
    .Y(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1031_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1796_  (.B1(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1037_ ),
    .VSS(VSS),
    .A1(net452),
    .A2(\i_ibex/ex_block_i/alu_i/_1030_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1797_  (.A(\i_ibex/ex_block_i/alu_i/_0687_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(net759),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1799_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/alu_operand_b_ex [22]),
    .A2(net601),
    .Y(\i_ibex/ex_block_i/alu_i/_1040_ ),
    .B1(net591));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_1800_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1041_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1040_ ),
    .A(net792));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1801_  (.A(\i_ibex/alu_operand_b_ex [22]),
    .B(net603),
    .Y(\i_ibex/ex_block_i/alu_i/_1042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1802_  (.B1(net804),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1043_ ),
    .VSS(VSS),
    .A1(net184),
    .A2(net185));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1803_  (.A(\i_ibex/ex_block_i/alu_i/_1042_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_1043_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1804_  (.A(net186),
    .B(net187),
    .X(\i_ibex/ex_block_i/alu_i/_1045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1805_  (.A(net579),
    .B(\i_ibex/alu_operand_b_ex [21]),
    .X(\i_ibex/ex_block_i/alu_i/_1046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1806_  (.A(net804),
    .B_N(net579),
    .Y(\i_ibex/ex_block_i/alu_i/_1047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1807_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net806),
    .A2(net188),
    .Y(\i_ibex/ex_block_i/alu_i/_1048_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1047_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1808_  (.A(\i_ibex/alu_operand_b_ex [21]),
    .B(net597),
    .C(\i_ibex/ex_block_i/alu_i/_1048_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1809_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1154),
    .C1(\i_ibex/ex_block_i/alu_i/_1049_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1046_ ),
    .A1(net791),
    .Y(\i_ibex/ex_block_i/alu_i/_1050_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1045_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1810_  (.A0(net591),
    .A1(net189),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_1051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1811_  (.B(net190),
    .C(net191),
    .A(net795),
    .Y(\i_ibex/ex_block_i/alu_i/_1052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1812_  (.B(\i_ibex/alu_operand_b_ex [22]),
    .C(net1154),
    .A(net592),
    .Y(\i_ibex/ex_block_i/alu_i/_1053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1813_  (.Y(\i_ibex/ex_block_i/alu_i/_1054_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1052_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1814_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1042_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1051_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1055_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1054_ ));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_1815_  (.Y(\i_ibex/ex_block_i/alu_i/_1056_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1050_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1055_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1044_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1816_  (.A2(\i_ibex/ex_block_i/alu_i/_1038_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1037_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1056_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1817_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_1057_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1058_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1023_ ),
    .A1(net981));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1818_  (.B1(\i_ibex/ex_block_i/alu_i/_1058_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1059_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0705_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1003_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1819_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/alu_operand_b_ex [26]),
    .A2(net602),
    .Y(\i_ibex/ex_block_i/alu_i/_1060_ ),
    .B1(net531));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1820_  (.B1(net805),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1061_ ),
    .VSS(VSS),
    .A1(net192),
    .A2(net193));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1821_  (.A(\i_ibex/ex_block_i/alu_i/_0635_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_1061_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1822_  (.B1(\i_ibex/ex_block_i/alu_i/_1062_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1063_ ),
    .VSS(VSS),
    .A1(net788),
    .A2(\i_ibex/ex_block_i/alu_i/_1060_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1823_  (.A0(net529),
    .A1(net194),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_1064_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1824_  (.A(net529),
    .B(\i_ibex/alu_operand_b_ex [25]),
    .X(\i_ibex/ex_block_i/alu_i/_1065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1825_  (.X(\i_ibex/ex_block_i/alu_i/_1066_ ),
    .A(net789),
    .B(net195),
    .C(net196),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1826_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1155),
    .C1(\i_ibex/ex_block_i/alu_i/_1066_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1065_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1064_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1067_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0643_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1827_  (.B(\i_ibex/alu_operand_b_ex [26]),
    .C(net1154),
    .A(net531),
    .Y(\i_ibex/ex_block_i/alu_i/_1068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1828_  (.A2(net601),
    .A1(\i_ibex/alu_operand_b_ex [25]),
    .B1(net529),
    .X(\i_ibex/ex_block_i/alu_i/_1069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1829_  (.B1(net793),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1070_ ),
    .VSS(VSS),
    .A1(net197),
    .A2(net198));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1830_  (.B1(\i_ibex/ex_block_i/alu_i/_1070_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1071_ ),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_b_ex [25]),
    .A2(net597));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1831_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1496),
    .A2(\i_ibex/ex_block_i/alu_i/_1069_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1072_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1071_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1832_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/alu_operand_b_ex [24]),
    .A2(net602),
    .Y(\i_ibex/ex_block_i/alu_i/_1073_ ),
    .B1(net527));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_1833_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1074_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1073_ ),
    .A(net795));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1834_  (.B1(net790),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1075_ ),
    .VSS(VSS),
    .A1(net199),
    .A2(net200));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1835_  (.A(\i_ibex/ex_block_i/alu_i/_0648_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_1075_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1836_  (.A0(net593),
    .A1(net201),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_1077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1837_  (.A(net593),
    .B(\i_ibex/alu_operand_b_ex [23]),
    .X(\i_ibex/ex_block_i/alu_i/_1078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1838_  (.X(\i_ibex/ex_block_i/alu_i/_1079_ ),
    .A(net800),
    .B(net202),
    .C(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1839_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1154),
    .C1(\i_ibex/ex_block_i/alu_i/_1079_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1078_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1077_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1080_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0656_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1840_  (.A0(net527),
    .A1(net204),
    .S(net788),
    .X(\i_ibex/ex_block_i/alu_i/_1081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1841_  (.A(net527),
    .B(\i_ibex/alu_operand_b_ex [24]),
    .X(\i_ibex/ex_block_i/alu_i/_1082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1842_  (.X(\i_ibex/ex_block_i/alu_i/_1083_ ),
    .A(net789),
    .B(net205),
    .C(net206),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1843_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1154),
    .C1(\i_ibex/ex_block_i/alu_i/_1083_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1082_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0648_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1084_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1081_ ));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_1844_  (.Y(\i_ibex/ex_block_i/alu_i/_1085_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1080_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1084_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1076_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1845_  (.Y(\i_ibex/ex_block_i/alu_i/_1086_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1085_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_1072_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1846_  (.A0(net531),
    .A1(net207),
    .S(net798),
    .X(\i_ibex/ex_block_i/alu_i/_1087_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1847_  (.A(net208),
    .B(net209),
    .X(\i_ibex/ex_block_i/alu_i/_1088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_1848_  (.Y(\i_ibex/ex_block_i/alu_i/_1089_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1088_ ),
    .B2(net792),
    .A2(\i_ibex/ex_block_i/alu_i/_1087_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0635_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_1849_  (.B(\i_ibex/ex_block_i/alu_i/_1068_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1086_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1067_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1090_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_1089_ ));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1850_  (.A(\i_ibex/ex_block_i/alu_i/_1063_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1090_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1091_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1851_  (.A2(\i_ibex/ex_block_i/alu_i/_1059_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0665_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1091_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout756 (.A(\i_ibex/id_stage_i/imm_u_type [22]),
    .X(net756),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net756),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(\i_ibex/id_stage_i/imm_u_type [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout753 (.A(\i_ibex/id_stage_i/imm_u_type [24]),
    .X(net753),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1856_  (.A(\i_ibex/alu_operand_b_ex [29]),
    .B(net604),
    .Y(\i_ibex/ex_block_i/alu_i/_1097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1857_  (.A(net210),
    .B(\i_ibex/ex_block_i/alu_i/_1097_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1858_  (.Y(\i_ibex/ex_block_i/alu_i/_1099_ ),
    .A(net211),
    .B(\i_ibex/ex_block_i/alu_i/_1098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(\i_ibex/id_stage_i/imm_u_type [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1860_  (.Y(\i_ibex/ex_block_i/alu_i/_1101_ ),
    .A(net560),
    .B(\i_ibex/alu_operand_b_ex [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1861_  (.Y(\i_ibex/ex_block_i/alu_i/_1102_ ),
    .A(net600),
    .B(\i_ibex/ex_block_i/alu_i/_1101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1862_  (.A(net802),
    .B(\i_ibex/ex_block_i/alu_i/_1102_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1863_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net808),
    .A2(\i_ibex/ex_block_i/alu_i/_1099_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1104_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1103_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1864_  (.A(\i_ibex/alu_operand_b_ex [30]),
    .B(net604),
    .Y(\i_ibex/ex_block_i/alu_i/_1105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1865_  (.A(net212),
    .B(\i_ibex/ex_block_i/alu_i/_1105_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1866_  (.Y(\i_ibex/ex_block_i/alu_i/_1107_ ),
    .A(net213),
    .B(\i_ibex/ex_block_i/alu_i/_1106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1867_  (.Y(\i_ibex/ex_block_i/alu_i/_1108_ ),
    .A(net581),
    .B(\i_ibex/alu_operand_b_ex [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1868_  (.Y(\i_ibex/ex_block_i/alu_i/_1109_ ),
    .A(net600),
    .B(\i_ibex/ex_block_i/alu_i/_1108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1869_  (.A(net802),
    .B(\i_ibex/ex_block_i/alu_i/_1109_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1870_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net808),
    .A2(\i_ibex/ex_block_i/alu_i/_1107_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1111_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1110_ ));
 sg13g2_buf_2 fanout751 (.A(net752),
    .X(net751),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1872_  (.Y(\i_ibex/ex_block_i/alu_i/_1113_ ),
    .A(net533),
    .B(\i_ibex/alu_operand_b_ex [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1873_  (.Y(\i_ibex/ex_block_i/alu_i/_1114_ ),
    .A(net599),
    .B(\i_ibex/ex_block_i/alu_i/_1113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1874_  (.A(\i_ibex/alu_operand_b_ex [27]),
    .B(net602),
    .Y(\i_ibex/ex_block_i/alu_i/_1115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1875_  (.A(net214),
    .B(\i_ibex/ex_block_i/alu_i/_1115_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1876_  (.Y(\i_ibex/ex_block_i/alu_i/_1117_ ),
    .A(net215),
    .B(\i_ibex/ex_block_i/alu_i/_1116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1877_  (.Y(\i_ibex/ex_block_i/alu_i/_1118_ ),
    .A(net806),
    .B(\i_ibex/ex_block_i/alu_i/_1117_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1878_  (.B1(\i_ibex/ex_block_i/alu_i/_1118_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .VSS(VSS),
    .A1(net801),
    .A2(\i_ibex/ex_block_i/alu_i/_1114_ ));
 sg13g2_buf_2 fanout750 (.A(net752),
    .X(net750),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1880_  (.Y(\i_ibex/ex_block_i/alu_i/_1121_ ),
    .A(net538),
    .B(\i_ibex/alu_operand_b_ex [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1881_  (.Y(\i_ibex/ex_block_i/alu_i/_1122_ ),
    .A(net599),
    .B(\i_ibex/ex_block_i/alu_i/_1121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1882_  (.A(\i_ibex/alu_operand_b_ex [28]),
    .B(net604),
    .Y(\i_ibex/ex_block_i/alu_i/_1123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1883_  (.A(net216),
    .B(\i_ibex/ex_block_i/alu_i/_1123_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1884_  (.Y(\i_ibex/ex_block_i/alu_i/_1125_ ),
    .A(net217),
    .B(\i_ibex/ex_block_i/alu_i/_1124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1885_  (.Y(\i_ibex/ex_block_i/alu_i/_1126_ ),
    .A(net807),
    .B(\i_ibex/ex_block_i/alu_i/_1125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1886_  (.B1(\i_ibex/ex_block_i/alu_i/_1126_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1127_ ),
    .VSS(VSS),
    .A1(net802),
    .A2(\i_ibex/ex_block_i/alu_i/_1122_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1887_  (.Y(\i_ibex/ex_block_i/alu_i/_1128_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1127_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1888_  (.A(\i_ibex/ex_block_i/alu_i/_1104_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1111_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1128_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1889_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/alu_operand_b_ex [28]),
    .C1(\i_ibex/ex_block_i/alu_i/_1123_ ),
    .B1(net1153),
    .A1(net806),
    .Y(\i_ibex/ex_block_i/alu_i/_1130_ ),
    .A2(net218));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1890_  (.A(net806),
    .B_N(net538),
    .Y(\i_ibex/ex_block_i/alu_i/_1131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1891_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net806),
    .A2(net219),
    .Y(\i_ibex/ex_block_i/alu_i/_1132_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1131_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1892_  (.A0(net533),
    .A1(net220),
    .S(net788),
    .X(\i_ibex/ex_block_i/alu_i/_1133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1893_  (.B(net221),
    .C(net222),
    .A(net806),
    .Y(\i_ibex/ex_block_i/alu_i/_1134_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1894_  (.B(\i_ibex/alu_operand_b_ex [27]),
    .C(net1153),
    .A(net533),
    .Y(\i_ibex/ex_block_i/alu_i/_1135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1895_  (.Y(\i_ibex/ex_block_i/alu_i/_1136_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1134_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1896_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1133_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1115_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1137_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1136_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1897_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1130_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1132_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1138_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1137_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1898_  (.A(\i_ibex/ex_block_i/alu_i/_1130_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1132_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1139_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1899_  (.A(\i_ibex/ex_block_i/alu_i/_1138_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1139_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1140_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout749 (.A(\i_ibex/id_stage_i/imm_u_type [26]),
    .X(net749),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1901_  (.A0(net561),
    .A1(net223),
    .S(net799),
    .X(\i_ibex/ex_block_i/alu_i/_1142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1902_  (.Y(\i_ibex/ex_block_i/alu_i/_1143_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1097_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1903_  (.B(net224),
    .C(net225),
    .A(net807),
    .Y(\i_ibex/ex_block_i/alu_i/_1144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1904_  (.B(\i_ibex/alu_operand_b_ex [29]),
    .C(net1153),
    .A(net561),
    .Y(\i_ibex/ex_block_i/alu_i/_1145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/ex_block_i/alu_i/_1905_  (.A(\i_ibex/ex_block_i/alu_i/_1140_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1143_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1144_ ),
    .D(\i_ibex/ex_block_i/alu_i/_1145_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1146_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1906_  (.A2(net601),
    .A1(\i_ibex/alu_operand_b_ex [29]),
    .B1(net561),
    .X(\i_ibex/ex_block_i/alu_i/_1147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1907_  (.B1(net807),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1148_ ),
    .VSS(VSS),
    .A1(net226),
    .A2(net227));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1908_  (.B1(\i_ibex/ex_block_i/alu_i/_1148_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1149_ ),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_b_ex [29]),
    .A2(net600));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1909_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1495),
    .A2(\i_ibex/ex_block_i/alu_i/_1147_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1150_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1149_ ));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net749),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1911_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/alu_operand_b_ex [30]),
    .A2(net604),
    .Y(\i_ibex/ex_block_i/alu_i/_1152_ ),
    .B1(net582));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1912_  (.B1(net807),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1153_ ),
    .VSS(VSS),
    .A1(net228),
    .A2(net229));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1913_  (.A(\i_ibex/ex_block_i/alu_i/_1105_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_1153_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1914_  (.B1(\i_ibex/ex_block_i/alu_i/_1154_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1155_ ),
    .VSS(VSS),
    .A1(net802),
    .A2(\i_ibex/ex_block_i/alu_i/_1152_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1915_  (.Y(\i_ibex/ex_block_i/alu_i/_1156_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1155_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_1150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1916_  (.A0(net582),
    .A1(net230),
    .S(net799),
    .X(\i_ibex/ex_block_i/alu_i/_1157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_1917_  (.A(net582),
    .B(\i_ibex/alu_operand_b_ex [30]),
    .X(\i_ibex/ex_block_i/alu_i/_1158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_1918_  (.X(\i_ibex/ex_block_i/alu_i/_1159_ ),
    .A(net802),
    .B(net231),
    .C(net232),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_1919_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_1158_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_1159_ ),
    .B1(net1153),
    .A1(\i_ibex/ex_block_i/alu_i/_1157_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1160_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1105_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1920_  (.B1(\i_ibex/ex_block_i/alu_i/_1160_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1161_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1146_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1156_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1921_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1092_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1129_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1162_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1161_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1922_  (.B(\i_ibex/alu_operand_b_ex [31]),
    .C(net600),
    .A(net1496),
    .Y(\i_ibex/ex_block_i/alu_i/_1163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1923_  (.B1(\i_ibex/ex_block_i/alu_i/_1163_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1164_ ),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_b_ex [31]),
    .A2(net600));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1924_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net808),
    .A2(net233),
    .Y(\i_ibex/ex_block_i/alu_i/_1165_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1164_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1925_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1166_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1165_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1926_  (.A0(net583),
    .A1(net234),
    .S(net799),
    .X(\i_ibex/ex_block_i/alu_i/_1167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1927_  (.A(\i_ibex/ex_block_i/alu_i/_1166_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1167_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1928_  (.Y(\i_ibex/ex_block_i/alu_i/_1169_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1166_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1929_  (.B1(\i_ibex/ex_block_i/alu_i/_1169_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_adder_result_ext [33]),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1162_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1168_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1930_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1170_ ),
    .A(net100),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1931_  (.Y(\i_ibex/ex_block_i/alu_i/_1171_ ),
    .A(net235),
    .B(net600),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1932_  (.B1(\i_ibex/ex_block_i/alu_i/_1171_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1172_ ),
    .VSS(VSS),
    .A1(net1495),
    .A2(net599));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1933_  (.B1(net808),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1173_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1170_ ),
    .A2(net236));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_1934_  (.Y(\i_ibex/ex_block_i/alu_i/_1174_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1173_ ),
    .B2(net604),
    .A2(\i_ibex/ex_block_i/alu_i/_1172_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1170_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1935_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_adder_result_ext [0]),
    .A(\i_ibex/ex_block_i/alu_i/_1174_ ),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_1936_  (.B(\i_ibex/ex_block_i/alu_i/_1167_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1165_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1937_  (.Y(\i_ibex/ex_block_i/alu_i/_1176_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1162_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/ex_block_i/alu_i/_1938_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [32]),
    .A(net1521),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1939_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1177_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0677_ ),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/ex_block_i/alu_i/_1940_  (.A(\i_ibex/ex_block_i/alu_i/_0901_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0969_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_1941_  (.A(\i_ibex/ex_block_i/alu_i/_1178_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_1002_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1179_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1942_  (.A(\i_ibex/ex_block_i/alu_i/_1021_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1179_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1180_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1943_  (.B1(\i_ibex/ex_block_i/alu_i/_1030_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1181_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0704_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1180_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1944_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1182_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1945_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1177_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1181_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1183_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1182_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1946_  (.B1(\i_ibex/ex_block_i/alu_i/_1050_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1184_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1183_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1947_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [23]),
    .A(\i_ibex/ex_block_i/alu_i/_0687_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_1948_  (.B(\i_ibex/ex_block_i/alu_i/_1183_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .X(\i_ibex/ex_block_i/alu_adder_result_ext [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1949_  (.A2(net601),
    .A1(\i_ibex/alu_operand_b_ex [19]),
    .B1(net575),
    .X(\i_ibex/ex_block_i/alu_i/_1185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1950_  (.B1(net791),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1186_ ),
    .VSS(VSS),
    .A1(net237),
    .A2(net238));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1951_  (.B1(\i_ibex/ex_block_i/alu_i/_1186_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1187_ ),
    .VSS(VSS),
    .A1(\i_ibex/alu_operand_b_ex [19]),
    .A2(net596));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1952_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_1187_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1185_ ),
    .A1(net1496));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1953_  (.Y(\i_ibex/ex_block_i/alu_i/_1189_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1003_ ),
    .A_N(net981),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_1954_  (.A0(\i_ibex/ex_block_i/alu_i/_1030_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .S(\i_ibex/ex_block_i/alu_i/_1189_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1955_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [21]),
    .A(\i_ibex/ex_block_i/alu_i/_1177_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1956_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [20]),
    .A(\i_ibex/ex_block_i/alu_i/_0704_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1957_  (.B1(\i_ibex/ex_block_i/alu_i/_1014_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1191_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1178_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0994_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1958_  (.Y(\i_ibex/ex_block_i/alu_i/_1192_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1959_  (.A(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1960_  (.A2(\i_ibex/ex_block_i/alu_i/_1192_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1191_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1193_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1961_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0985_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1194_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1195_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1009_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1962_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [19]),
    .A(\i_ibex/ex_block_i/alu_i/_0977_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1195_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1963_  (.B1(\i_ibex/ex_block_i/alu_i/_1192_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1196_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1191_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1193_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1964_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [18]),
    .A(\i_ibex/ex_block_i/alu_i/_0985_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1965_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [17]),
    .A(\i_ibex/ex_block_i/alu_i/_1001_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1191_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1966_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1197_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0994_ ),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1967_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [16]),
    .A(\i_ibex/ex_block_i/alu_i/_1178_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1968_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1198_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0932_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1969_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1199_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_1970_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1200_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0849_ ),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/ex_block_i/alu_i/_1971_  (.A(\i_ibex/ex_block_i/alu_i/_0713_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0717_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1201_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1972_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0744_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0841_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1202_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1201_ ));
 sg13g2_a21oi_2 \i_ibex/ex_block_i/alu_i/_1973_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/ex_block_i/alu_i/_0963_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1203_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1202_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1200_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1974_  (.B1(\i_ibex/ex_block_i/alu_i/_0943_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1204_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1199_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1203_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_1975_  (.B(\i_ibex/ex_block_i/alu_i/_0946_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0948_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0945_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1976_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0857_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1204_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1206_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1205_ ));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_1977_  (.A(\i_ibex/ex_block_i/alu_i/_0881_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0898_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1206_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1978_  (.A(\i_ibex/ex_block_i/alu_i/_1198_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1207_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1208_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1979_  (.B1(\i_ibex/ex_block_i/alu_i/_0934_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1209_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1208_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1980_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [15]),
    .A(\i_ibex/ex_block_i/alu_i/_0873_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_1981_  (.B(\i_ibex/ex_block_i/alu_i/_1208_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .X(\i_ibex/ex_block_i/alu_adder_result_ext [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1982_  (.Y(\i_ibex/ex_block_i/alu_i/_1210_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0665_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_1983_  (.A2(\i_ibex/ex_block_i/alu_i/_1023_ ),
    .A1(net981),
    .B1(\i_ibex/ex_block_i/alu_i/_1057_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1984_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0665_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1211_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1212_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1091_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1985_  (.B1(\i_ibex/ex_block_i/alu_i/_1212_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1213_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1003_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1210_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1986_  (.Y(\i_ibex/ex_block_i/alu_i/_1214_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1213_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_1128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_1987_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1146_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1214_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1215_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1150_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1988_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [31]),
    .A(\i_ibex/ex_block_i/alu_i/_1111_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1215_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_1989_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1216_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1206_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0881_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_1990_  (.Y(\i_ibex/ex_block_i/alu_i/_1217_ ),
    .B(net1158),
    .A_N(\i_ibex/ex_block_i/alu_i/_0922_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_1991_  (.B1(\i_ibex/ex_block_i/alu_i/_1217_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1218_ ),
    .VSS(VSS),
    .A1(net1158),
    .A2(\i_ibex/ex_block_i/alu_i/_0910_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1992_  (.Y(\i_ibex/ex_block_i/alu_i/_1219_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1216_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1218_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1993_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [13]),
    .A(\i_ibex/ex_block_i/alu_i/_0898_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1219_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_1994_  (.Y(\i_ibex/ex_block_i/alu_i/_1220_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0857_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_1995_  (.A(\i_ibex/ex_block_i/alu_i/_1220_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1203_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1221_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_1996_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1222_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1221_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0950_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1997_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [12]),
    .A(\i_ibex/ex_block_i/alu_i/_0881_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1222_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1998_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [11]),
    .A(\i_ibex/ex_block_i/alu_i/_0936_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_1999_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [10]),
    .A(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2000_  (.Y(\i_ibex/ex_block_i/alu_i/_1223_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0954_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_1202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2001_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [9]),
    .A(\i_ibex/ex_block_i/alu_i/_0849_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2002_  (.Y(\i_ibex/ex_block_i/alu_i/_1224_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0744_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0841_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2003_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [8]),
    .A(\i_ibex/ex_block_i/alu_i/_1201_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1224_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2004_  (.Y(\i_ibex/ex_block_i/alu_i/_1225_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0824_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0840_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2005_  (.B1(\i_ibex/ex_block_i/alu_i/_0727_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1226_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0751_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1225_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2006_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [7]),
    .A(\i_ibex/ex_block_i/alu_i/_0757_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1226_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2007_  (.A2(\i_ibex/ex_block_i/alu_i/_0747_ ),
    .A1(net807),
    .B1(\i_ibex/ex_block_i/alu_i/_0750_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2008_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [6]),
    .A(\i_ibex/ex_block_i/alu_i/_1227_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/ex_block_i/alu_i/_2009_  (.Y(\i_ibex/ex_block_i/alu_i/_1228_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0782_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0823_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2010_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1229_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0838_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0835_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2011_  (.A2(\i_ibex/ex_block_i/alu_i/_1229_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1228_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0832_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1230_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2012_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [5]),
    .A(\i_ibex/ex_block_i/alu_i/_0831_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1230_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2013_  (.B(\i_ibex/ex_block_i/alu_i/_1229_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1228_ ),
    .X(\i_ibex/ex_block_i/alu_adder_result_ext [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2014_  (.Y(\i_ibex/ex_block_i/alu_i/_1231_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1140_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1214_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2015_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [30]),
    .A(\i_ibex/ex_block_i/alu_i/_1104_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2016_  (.A(\i_ibex/ex_block_i/alu_i/_0785_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0788_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1232_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2017_  (.B(net526),
    .A(net536),
    .X(\i_ibex/ex_block_i/alu_i/_1233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2018_  (.A0(net239),
    .A1(\i_ibex/ex_block_i/alu_i/_1233_ ),
    .S(net1495),
    .X(\i_ibex/ex_block_i/alu_i/_1234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2019_  (.Y(\i_ibex/ex_block_i/alu_i/_1235_ ),
    .A(net791),
    .B(net526),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2020_  (.Y(\i_ibex/ex_block_i/alu_i/_1236_ ),
    .B1(net1158),
    .B2(\i_ibex/ex_block_i/alu_i/_1235_ ),
    .A2(net240),
    .A1(net803),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2021_  (.B(\i_ibex/ex_block_i/alu_i/_1236_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1234_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/ex_block_i/alu_i/_2022_  (.Y(\i_ibex/ex_block_i/alu_i/_1238_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0801_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0803_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2023_  (.A(net599),
    .B(\i_ibex/ex_block_i/alu_i/_1238_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1239_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2024_  (.A(\i_ibex/ex_block_i/alu_i/_0809_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1239_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1240_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2025_  (.Y(\i_ibex/ex_block_i/alu_i/_1241_ ),
    .A(net1157),
    .B(\i_ibex/ex_block_i/alu_i/_0813_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2026_  (.B1(\i_ibex/ex_block_i/alu_i/_1241_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1242_ ),
    .VSS(VSS),
    .A1(net1157),
    .A2(\i_ibex/ex_block_i/alu_i/_0819_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2027_  (.B1(\i_ibex/ex_block_i/alu_i/_1242_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1243_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1237_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1240_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2028_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [3]),
    .A(\i_ibex/ex_block_i/alu_i/_1232_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1243_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2029_  (.A(net241),
    .B(\i_ibex/ex_block_i/alu_i/_1235_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2030_  (.Y(\i_ibex/ex_block_i/alu_i/_1245_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1238_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2031_  (.Y(\i_ibex/ex_block_i/alu_i/_1246_ ),
    .A(net805),
    .B(net242),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2032_  (.Y(\i_ibex/ex_block_i/alu_i/_1247_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0809_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2033_  (.Y(\i_ibex/ex_block_i/alu_i/_1248_ ),
    .A(net603),
    .B(\i_ibex/ex_block_i/alu_i/_1247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2034_  (.B1(\i_ibex/ex_block_i/alu_i/_1248_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1249_ ),
    .VSS(VSS),
    .A1(net599),
    .A2(\i_ibex/ex_block_i/alu_i/_1245_ ));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2035_  (.B(\i_ibex/ex_block_i/alu_i/_1249_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1234_ ),
    .X(\i_ibex/ex_block_i/alu_adder_result_ext [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2036_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1052),
    .A2(net1157),
    .Y(\i_ibex/ex_block_i/alu_i/_1250_ ),
    .B1(net243));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2037_  (.Y(\i_ibex/ex_block_i/alu_i/_1251_ ),
    .A(net100),
    .B(net244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2038_  (.Y(\i_ibex/ex_block_i/alu_i/_1252_ ),
    .B(net245),
    .A_N(net246),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2039_  (.B1(\i_ibex/ex_block_i/alu_i/_1252_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1253_ ),
    .VSS(VSS),
    .A1(net247),
    .A2(\i_ibex/ex_block_i/alu_i/_1251_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2040_  (.Y(\i_ibex/ex_block_i/alu_i/_1254_ ),
    .A(net602),
    .B(\i_ibex/ex_block_i/alu_i/_1253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2041_  (.B1(\i_ibex/ex_block_i/alu_i/_1254_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1255_ ),
    .VSS(VSS),
    .A1(net100),
    .A2(\i_ibex/ex_block_i/alu_i/_1250_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2042_  (.Y(\i_ibex/ex_block_i/alu_i/_1256_ ),
    .B(net100),
    .A_N(net248),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2043_  (.B1(net792),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1257_ ),
    .VSS(VSS),
    .A1(net599),
    .A2(\i_ibex/ex_block_i/alu_i/_1256_ ));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2044_  (.Y(\i_ibex/ex_block_i/alu_i/_1258_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1257_ ),
    .B2(net488),
    .A2(\i_ibex/ex_block_i/alu_i/_1255_ ),
    .A1(net803),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2045_  (.A0(net535),
    .A1(net249),
    .S(net787),
    .X(\i_ibex/ex_block_i/alu_i/_1259_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2046_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [1]),
    .A(\i_ibex/ex_block_i/alu_i/_1258_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1259_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2047_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_1213_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_1136_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1133_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1260_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1115_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2048_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [29]),
    .A(\i_ibex/ex_block_i/alu_i/_1127_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2049_  (.B(\i_ibex/ex_block_i/alu_i/_1213_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .X(\i_ibex/ex_block_i/alu_adder_result_ext [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2050_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0664_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1059_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1261_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1085_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2051_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1067_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1261_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1262_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1072_ ));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2052_  (.B(\i_ibex/ex_block_i/alu_i/_1262_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0639_ ),
    .X(\i_ibex/ex_block_i/alu_adder_result_ext [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2053_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [26]),
    .A(\i_ibex/ex_block_i/alu_i/_0647_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2054_  (.Y(\i_ibex/ex_block_i/alu_i/_1263_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1059_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_0663_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2055_  (.Y(\i_ibex/ex_block_i/alu_i/_1264_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1080_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1263_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2056_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [25]),
    .A(\i_ibex/ex_block_i/alu_i/_0655_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2057_  (.Y(\i_ibex/ex_block_i/alu_adder_result_ext [24]),
    .A(\i_ibex/ex_block_i/alu_i/_0663_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout747 (.A(net749),
    .X(net747),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/ex_block_i/alu_i/_2059_  (.A(\i_ibex/alu_operand_b_ex [31]),
    .B_N(net583),
    .Y(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2060_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1267_ ),
    .A(net1292),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2061_  (.A(net325),
    .B(\i_ibex/alu_operator_ex [4]),
    .Y(\i_ibex/ex_block_i/alu_i/_1268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2062_  (.A(\i_ibex/alu_operator_ex [5]),
    .B(\i_ibex/ex_block_i/alu_i/_1268_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1269_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/ex_block_i/alu_i/_2063_  (.Y(\i_ibex/ex_block_i/alu_i/_1270_ ),
    .A(net622),
    .B(\i_ibex/ex_block_i/alu_i/_0597_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2064_  (.Y(\i_ibex/ex_block_i/alu_i/_1271_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_0605_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2065_  (.B1(\i_ibex/ex_block_i/alu_i/_1271_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1272_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1270_ ));
 sg13g2_nor2_2 \i_ibex/ex_block_i/alu_i/_2066_  (.A(net326),
    .B(\i_ibex/ex_block_i/alu_i/_0612_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1273_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(\i_ibex/id_stage_i/imm_u_type [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2068_  (.B(\i_ibex/ex_block_i/alu_i/_1270_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0605_ ),
    .A(net1289),
    .Y(\i_ibex/ex_block_i/alu_i/_1275_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2069_  (.B1(\i_ibex/ex_block_i/alu_i/_1275_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1276_ ),
    .VSS(VSS),
    .A1(net1289),
    .A2(\i_ibex/ex_block_i/alu_i/_1270_ ));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2070_  (.Y(\i_ibex/ex_block_i/alu_i/_1277_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1273_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1276_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1272_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1269_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2071_  (.A(net622),
    .B(net1290),
    .Y(\i_ibex/ex_block_i/alu_i/_1278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2072_  (.A(\i_ibex/ex_block_i/alu_i/_1267_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1269_ ),
    .X(\i_ibex/ex_block_i/alu_i/_1279_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2073_  (.B(\i_ibex/ex_block_i/alu_i/_1278_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1279_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1280_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2074_  (.B1(\i_ibex/ex_block_i/alu_i/_1280_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1281_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1267_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1277_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2075_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1282_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1281_ ),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2076_  (.Y(\i_ibex/ex_block_i/alu_i/_1283_ ),
    .A(net622),
    .B(net1292),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2077_  (.Y(\i_ibex/ex_block_i/alu_i/_1284_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1283_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1269_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1273_ ),
    .A1(net1292),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2078_  (.A(net1290),
    .B(\i_ibex/ex_block_i/alu_i/_1284_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1285_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_2079_  (.X(\i_ibex/ex_block_i/alu_i/_1286_ ),
    .A(net621),
    .B(net1293),
    .C(\i_ibex/ex_block_i/alu_i/_1273_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2080_  (.B1(net1289),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1287_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1285_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1286_ ));
 sg13g2_buf_2 fanout745 (.A(net746),
    .X(net745),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2082_  (.Y(\i_ibex/ex_block_i/alu_i/_1289_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1282_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1287_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2083_  (.Y(\i_ibex/ex_block_i/alu_i/_1290_ ),
    .A(net1288),
    .B(net622),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2084_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1291_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1290_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2085_  (.Y(\i_ibex/ex_block_i/alu_i/_1292_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1291_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1279_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1286_ ),
    .A1(net1288),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2086_  (.A(net1289),
    .B(net621),
    .Y(\i_ibex/ex_block_i/alu_i/_1293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_2087_  (.B(net1292),
    .C(\i_ibex/ex_block_i/alu_i/_1273_ ),
    .A(net1291),
    .Y(\i_ibex/ex_block_i/alu_i/_1294_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_1293_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2088_  (.B1(\i_ibex/ex_block_i/alu_i/_1294_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1295_ ),
    .VSS(VSS),
    .A1(net1290),
    .A2(\i_ibex/ex_block_i/alu_i/_1292_ ));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2089_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1296_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1295_ ),
    .A(net1151));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2090_  (.A0(\i_ibex/ex_block_i/alu_i/_1289_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1296_ ),
    .S(net1522),
    .X(\i_ibex/ex_block_i/alu_i/_1297_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2091_  (.A(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1297_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1298_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2092_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1299_ ),
    .A(\i_ibex/alu_operand_b_ex [31]),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/ex_block_i/alu_i/_2093_  (.A(net583),
    .B(\i_ibex/ex_block_i/alu_i/_1299_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2094_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_1301_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1287_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1281_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2095_  (.A(net1290),
    .B(\i_ibex/ex_block_i/alu_i/_1292_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/ex_block_i/alu_i/_2096_  (.A(\i_ibex/ex_block_i/alu_i/_1302_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_1294_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2097_  (.Y(\i_ibex/ex_block_i/alu_i/_1304_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1287_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2098_  (.A0(\i_ibex/ex_block_i/alu_i/_1301_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1304_ ),
    .S(net1522),
    .X(\i_ibex/ex_block_i/alu_i/_1305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2099_  (.A0(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .S(net1151),
    .X(\i_ibex/ex_block_i/alu_i/_1306_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2100_  (.A0(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .S(net1151),
    .X(\i_ibex/ex_block_i/alu_i/_1307_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2101_  (.Y(\i_ibex/ex_block_i/alu_i/_1308_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1307_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1282_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1306_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2102_  (.B1(\i_ibex/ex_block_i/alu_i/_1308_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1309_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1305_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2103_  (.Y(\i_ibex/ex_block_i/alu_i/_1310_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0603_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0615_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2104_  (.A(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1311_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2105_  (.A(\i_ibex/ex_block_i/alu_i/_1299_ ),
    .B(net1151),
    .X(\i_ibex/ex_block_i/alu_i/_1312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2106_  (.A(net583),
    .B(\i_ibex/ex_block_i/alu_i/_1299_ ),
    .C(net1151),
    .Y(\i_ibex/ex_block_i/alu_i/_1313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2107_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net583),
    .C1(\i_ibex/ex_block_i/alu_i/_1313_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1312_ ),
    .A1(net1521),
    .Y(\i_ibex/ex_block_i/alu_i/_1314_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1311_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2108_  (.Y(\i_ibex/ex_block_i/alu_i/_1315_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1281_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2109_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net584),
    .A2(\i_ibex/ex_block_i/alu_i/_1312_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1316_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1313_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2110_  (.Y(\i_ibex/ex_block_i/alu_i/_1317_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1295_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1316_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2111_  (.B1(\i_ibex/ex_block_i/alu_i/_1317_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1318_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1295_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1310_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2112_  (.A(\i_ibex/ex_block_i/alu_i/_1303_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1307_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2113_  (.Y(\i_ibex/ex_block_i/alu_i/_1320_ ),
    .A(net1521),
    .B(\i_ibex/ex_block_i/alu_i/_1319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2114_  (.B(\i_ibex/ex_block_i/alu_i/_1318_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1320_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1282_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2115_  (.B1(\i_ibex/ex_block_i/alu_i/_1321_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1322_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1314_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1315_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2116_  (.B(\i_ibex/ex_block_i/alu_i/_1198_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1218_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0898_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2117_  (.Y(\i_ibex/ex_block_i/alu_i/_1324_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0898_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1218_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2118_  (.B(\i_ibex/ex_block_i/alu_i/_0932_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1324_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1325_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2119_  (.B1(\i_ibex/ex_block_i/alu_i/_1325_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1326_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1323_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2120_  (.B1(\i_ibex/ex_block_i/alu_i/_1216_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1327_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0932_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1218_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2121_  (.A(\i_ibex/ex_block_i/alu_i/_0889_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0898_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1328_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2122_  (.Y(\i_ibex/ex_block_i/alu_i/_1329_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1327_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1328_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1326_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2123_  (.B(\i_ibex/ex_block_i/alu_i/_0647_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0664_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0639_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2124_  (.Y(\i_ibex/ex_block_i/alu_i/_1331_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1091_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2125_  (.A(\i_ibex/ex_block_i/alu_i/_0705_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1003_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1332_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2126_  (.Y(\i_ibex/ex_block_i/alu_i/_1333_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0665_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1332_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2127_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1331_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1333_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1334_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1119_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2128_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1335_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1178_ ),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2129_  (.A(\i_ibex/ex_block_i/alu_i/_1009_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1192_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2130_  (.Y(\i_ibex/ex_block_i/alu_i/_1337_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0977_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2131_  (.Y(\i_ibex/ex_block_i/alu_i/_1338_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0985_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_1014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2132_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1339_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0985_ ),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2133_  (.B(\i_ibex/ex_block_i/alu_i/_1014_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1339_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1340_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2134_  (.B1(\i_ibex/ex_block_i/alu_i/_1340_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_1341_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1338_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2135_  (.Y(\i_ibex/ex_block_i/alu_i/_1342_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0997_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2136_  (.A(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1339_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1342_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2137_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1000_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1341_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1344_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1343_ ));
 sg13g2_nor4_1 \i_ibex/ex_block_i/alu_i/_2138_  (.A(\i_ibex/ex_block_i/alu_i/_1335_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1197_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1337_ ),
    .D(\i_ibex/ex_block_i/alu_i/_1344_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1345_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2139_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net981),
    .A2(\i_ibex/ex_block_i/alu_i/_1345_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_1346_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1179_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2140_  (.Y(\i_ibex/ex_block_i/alu_i/_1347_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1345_ ),
    .A_N(net981),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2141_  (.A0(\i_ibex/ex_block_i/alu_i/_1346_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1347_ ),
    .S(\i_ibex/ex_block_i/alu_i/_0704_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2142_  (.Y(\i_ibex/ex_block_i/alu_i/_0001_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0677_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2143_  (.B(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .A(net452),
    .X(\i_ibex/ex_block_i/alu_i/_0002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2144_  (.A(\i_ibex/ex_block_i/alu_i/_1030_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0704_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2145_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0004_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0003_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0677_ ));
 sg13g2_a22oi_1 \i_ibex/ex_block_i/alu_i/_2146_  (.Y(\i_ibex/ex_block_i/alu_i/_0005_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0004_ ),
    .B2(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0002_ ),
    .A1(net981),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2147_  (.B1(\i_ibex/ex_block_i/alu_i/_0005_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0006_ ),
    .VSS(VSS),
    .A1(net981),
    .A2(\i_ibex/ex_block_i/alu_i/_0001_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2148_  (.Y(\i_ibex/ex_block_i/alu_i/_0007_ ),
    .A(net452),
    .B(\i_ibex/ex_block_i/alu_i/_1030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2149_  (.A(net452),
    .B(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2150_  (.A(net452),
    .B(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2151_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0003_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0008_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0010_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0009_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2152_  (.A0(\i_ibex/ex_block_i/alu_i/_0007_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0010_ ),
    .S(net981),
    .X(\i_ibex/ex_block_i/alu_i/_0011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_2153_  (.B(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0012_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/ex_block_i/alu_i/_0011_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2154_  (.B1(\i_ibex/ex_block_i/alu_i/_0012_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0013_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0006_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2155_  (.Y(\i_ibex/ex_block_i/alu_i/_0014_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2156_  (.B(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0014_ ),
    .A(net452),
    .Y(\i_ibex/ex_block_i/alu_i/_0015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2157_  (.Y(\i_ibex/ex_block_i/alu_i/_0016_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1036_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2158_  (.Y(\i_ibex/ex_block_i/alu_i/_0017_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0695_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_2159_  (.A(net452),
    .B(\i_ibex/ex_block_i/alu_i/_1188_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0017_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2160_  (.B(\i_ibex/ex_block_i/alu_i/_0015_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0018_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1179_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2161_  (.B1(\i_ibex/ex_block_i/alu_i/_0019_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0020_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1179_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0013_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2162_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0021_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0664_ ),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2163_  (.Y(\i_ibex/ex_block_i/alu_i/_0022_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1080_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0655_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_2164_  (.B(\i_ibex/ex_block_i/alu_i/_0663_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1058_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1091_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0023_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0022_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2165_  (.B1(\i_ibex/ex_block_i/alu_i/_0023_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0024_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0021_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1058_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2166_  (.Y(\i_ibex/ex_block_i/alu_i/_0025_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0663_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2167_  (.A(\i_ibex/ex_block_i/alu_i/_1091_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0025_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2168_  (.A(\i_ibex/ex_block_i/alu_i/_0021_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0665_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1058_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2169_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_1058_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0027_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0026_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0028_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0024_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2170_  (.A0(\i_ibex/ex_block_i/alu_i/_0028_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0021_ ),
    .S(\i_ibex/ex_block_i/alu_i/_1332_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2171_  (.Y(\i_ibex/ex_block_i/alu_i/_0030_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0849_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2172_  (.A(\i_ibex/ex_block_i/alu_i/_1201_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_0758_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2173_  (.Y(\i_ibex/ex_block_i/alu_i/_0032_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1201_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0743_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2174_  (.B(\i_ibex/ex_block_i/alu_i/_0757_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0032_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0727_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2175_  (.Y(\i_ibex/ex_block_i/alu_i/_0034_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0743_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0736_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2176_  (.Y(\i_ibex/ex_block_i/alu_i/_0035_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1201_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_2177_  (.A(\i_ibex/ex_block_i/alu_i/_0727_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0757_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0035_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2178_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0033_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0036_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0037_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1227_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2179_  (.A0(\i_ibex/ex_block_i/alu_i/_0031_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0037_ ),
    .S(\i_ibex/ex_block_i/alu_i/_1225_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_2180_  (.B(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0958_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0039_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/ex_block_i/alu_i/_1223_ ));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2181_  (.Y(\i_ibex/ex_block_i/alu_i/_0040_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0832_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0831_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_2182_  (.A(\i_ibex/ex_block_i/alu_i/_1228_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1229_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0040_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2183_  (.A2(\i_ibex/ex_block_i/alu_i/_0827_ ),
    .A1(net807),
    .B1(\i_ibex/ex_block_i/alu_i/_0830_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2184_  (.B(\i_ibex/ex_block_i/alu_i/_0042_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1229_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1228_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_2185_  (.B(\i_ibex/ex_block_i/alu_i/_1330_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1119_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0044_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/ex_block_i/alu_i/_1091_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2186_  (.A(\i_ibex/ex_block_i/alu_i/_0857_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1205_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2187_  (.Y(\i_ibex/ex_block_i/alu_i/_0046_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0881_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2188_  (.A(net1157),
    .B(\i_ibex/ex_block_i/alu_i/_0819_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0809_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2189_  (.B(\i_ibex/ex_block_i/alu_i/_0813_ ),
    .C(\i_ibex/ex_block_i/alu_i/_1238_ ),
    .A(net1157),
    .Y(\i_ibex/ex_block_i/alu_i/_0048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2190_  (.A(\i_ibex/ex_block_i/alu_i/_0047_ ),
    .B_N(\i_ibex/ex_block_i/alu_i/_0048_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2191_  (.Y(\i_ibex/ex_block_i/alu_i/_0050_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1232_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2192_  (.A(\i_ibex/ex_block_i/alu_i/_0864_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0962_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/ex_block_i/alu_i/_2193_  (.A(net435),
    .B(\i_ibex/ex_block_i/alu_adder_result_ext [1]),
    .C(\i_ibex/ex_block_i/alu_i/_0050_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0051_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2194_  (.B(\i_ibex/ex_block_i/alu_i/_0046_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0052_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0044_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2195_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0041_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0043_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0054_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0053_ ));
 sg13g2_nand4_1 \i_ibex/ex_block_i/alu_i/_2196_  (.B(\i_ibex/ex_block_i/alu_i/_0038_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0039_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0030_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0055_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0054_ ));
 sg13g2_or4_1 \i_ibex/ex_block_i/alu_i/_2197_  (.A(\i_ibex/ex_block_i/alu_adder_result_ext [11]),
    .B(\i_ibex/ex_block_i/alu_i/_0020_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0029_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0055_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/ex_block_i/alu_i/_2198_  (.A(\i_ibex/ex_block_i/alu_adder_result_ext [30]),
    .B(\i_ibex/ex_block_i/alu_i/_1334_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0000_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0056_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2199_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0058_ ),
    .B(\i_ibex/ex_block_i/alu_adder_result_ext [26]),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [29]));
 sg13g2_or4_1 \i_ibex/ex_block_i/alu_i/_2200_  (.A(\i_ibex/ex_block_i/alu_adder_result_ext [31]),
    .B(\i_ibex/ex_block_i/alu_i/_1329_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0057_ ),
    .D(\i_ibex/ex_block_i/alu_i/_0058_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2201_  (.Y(\i_ibex/ex_block_i/alu_i/_0060_ ),
    .B(net1521),
    .A_N(\i_ibex/ex_block_i/alu_adder_result_ext [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/ex_block_i/alu_i/_2202_  (.A(\i_ibex/ex_block_i/alu_adder_result_ext [23]),
    .B(\i_ibex/ex_block_i/alu_adder_result_ext [15]),
    .C(\i_ibex/ex_block_i/alu_i/_0059_ ),
    .Y(\i_ibex/ex_block_i/alu_is_equal_result ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0060_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2203_  (.A0(\i_ibex/ex_block_i/alu_i/_1310_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1322_ ),
    .S(\i_ibex/ex_block_i/alu_is_equal_result ),
    .X(\i_ibex/ex_block_i/alu_i/_0061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2204_  (.B1(\i_ibex/ex_block_i/alu_i/_0061_ ),
    .VDD(VDD),
    .Y(\i_ibex/branch_decision ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_1298_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1309_ ));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2205_  (.B(net1292),
    .C(\i_ibex/ex_block_i/alu_i/_1293_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0597_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2206_  (.B1(\i_ibex/ex_block_i/alu_i/_0062_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0063_ ),
    .VSS(VSS),
    .A1(net1292),
    .A2(\i_ibex/ex_block_i/alu_i/_0614_ ));
 sg13g2_nor4_2 \i_ibex/ex_block_i/alu_i/_2207_  (.A(net327),
    .B(\i_ibex/alu_operator_ex [4]),
    .C(\i_ibex/alu_operator_ex [5]),
    .Y(\i_ibex/ex_block_i/alu_i/_0064_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net1292));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2208_  (.A(\i_ibex/ex_block_i/alu_i/_1278_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0064_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2209_  (.A2(\i_ibex/ex_block_i/alu_i/_0063_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1273_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0065_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0066_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2210_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0067_ ),
    .B(net621),
    .A(net1288));
 sg13g2_nand3b_1 \i_ibex/ex_block_i/alu_i/_2211_  (.B(net1292),
    .C(\i_ibex/ex_block_i/alu_i/_1268_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/alu_operator_ex [5]));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2212_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1290),
    .A2(\i_ibex/ex_block_i/alu_i/_0067_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0069_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0068_ ));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2213_  (.Y(\i_ibex/ex_block_i/alu_i/_0070_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0064_ ),
    .A_N(\i_ibex/ex_block_i/alu_i/_1278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/ex_block_i/alu_i/_2214_  (.Y(\i_ibex/ex_block_i/alu_i/_0071_ ),
    .A(net1213),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/ex_block_i/alu_i/_2215_  (.A(\i_ibex/ex_block_i/alu_i/_0611_ ),
    .B(net1149),
    .C(net1180),
    .Y(\i_ibex/ex_block_i/alu_i/_0072_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/ex_block_i/alu_i/_0071_ ));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(\i_ibex/id_stage_i/imm_u_type [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout743 (.A(\i_ibex/id_stage_i/imm_u_type [28]),
    .X(net743),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(\i_ibex/id_stage_i/imm_u_type [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/ex_block_i/alu_i/_2219_  (.A(net1288),
    .B(\i_ibex/ex_block_i/alu_i/_1270_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0068_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout741 (.A(net742),
    .X(net741),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout740 (.A(\i_ibex/instr_rdata_id [2]),
    .X(net740),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout738 (.A(net740),
    .X(net738),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2224_  (.A(\i_ibex/alu_operand_b_ex [2]),
    .B(net526),
    .C(net489),
    .Y(\i_ibex/ex_block_i/alu_i/_0081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2225_  (.A(net697),
    .B(\i_ibex/ex_block_i/alu_i/_0081_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2226_  (.Y(\i_ibex/ex_block_i/alu_i/_0083_ ),
    .A(\i_ibex/alu_operand_b_ex [3]),
    .B(\i_ibex/ex_block_i/alu_i/_0082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout737 (.A(\i_ibex/id_stage_i/imm_u_type [30]),
    .X(net737),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2228_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0085_ ),
    .A(\i_ibex/alu_operand_b_ex [3]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2229_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0085_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0081_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0086_ ),
    .B1(net697));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2230_  (.Y(\i_ibex/ex_block_i/alu_i/_0087_ ),
    .A(\i_ibex/alu_operand_b_ex [4]),
    .B(\i_ibex/ex_block_i/alu_i/_0086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2231_  (.A(net439),
    .B(net996),
    .X(\i_ibex/ex_block_i/alu_i/_0088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2232_  (.A(net1288),
    .B(\i_ibex/ex_block_i/alu_i/_1270_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0068_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0089_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2233_  (.A0(net583),
    .A1(net535),
    .S(net1203),
    .X(\i_ibex/ex_block_i/alu_i/_0090_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/ex_block_i/alu_i/_2234_  (.A(net1290),
    .B(\i_ibex/ex_block_i/alu_i/_0067_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0068_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0091_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout736 (.A(net737),
    .X(net736),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2236_  (.A(net1052),
    .B(net697),
    .Y(\i_ibex/ex_block_i/alu_i/_0093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2237_  (.Y(\i_ibex/ex_block_i/alu_i/_0094_ ),
    .A(net526),
    .B(\i_ibex/ex_block_i/alu_i/_0093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout735 (.A(net737),
    .X(net735),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2239_  (.A(net526),
    .B(net488),
    .Y(\i_ibex/ex_block_i/alu_i/_0096_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2240_  (.A(net697),
    .B(\i_ibex/ex_block_i/alu_i/_0096_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2241_  (.Y(\i_ibex/ex_block_i/alu_i/_0098_ ),
    .A(\i_ibex/alu_operand_b_ex [2]),
    .B(\i_ibex/ex_block_i/alu_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2242_  (.Y(\i_ibex/ex_block_i/alu_i/_0099_ ),
    .A(net1017),
    .B(net1011),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2243_  (.A(net488),
    .B(\i_ibex/ex_block_i/alu_i/_0099_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0100_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2244_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0101_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0100_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0091_ ));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2245_  (.A(\i_ibex/ex_block_i/alu_i/_0090_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0101_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/ex_block_i/alu_i/_2246_  (.A(\i_ibex/ex_block_i/alu_i/_0090_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0091_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2247_  (.A(\i_ibex/ex_block_i/alu_i/_0088_ ),
    .B_N(net1087),
    .Y(\i_ibex/ex_block_i/alu_i/_0104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2248_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0088_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0102_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0105_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0104_ ));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(net737),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout733 (.A(\i_ibex/id_stage_i/imm_u_type [31]),
    .X(net733),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout732 (.A(net733),
    .X(net732),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net732),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2253_  (.S0(net1050),
    .A0(net550),
    .A1(net548),
    .A2(net527),
    .A3(net530),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2254_  (.S0(net1209),
    .A0(net560),
    .A1(net540),
    .A2(net538),
    .A3(net543),
    .S1(net490),
    .X(\i_ibex/ex_block_i/alu_i/_0111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2255_  (.S0(net1051),
    .A0(net546),
    .A1(net544),
    .A2(net531),
    .A3(net534),
    .S1(net1199),
    .X(\i_ibex/ex_block_i/alu_i/_0112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2256_  (.S0(net487),
    .A0(net585),
    .A1(net581),
    .A2(net535),
    .A3(net537),
    .S1(net1209),
    .X(\i_ibex/ex_block_i/alu_i/_0113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout730 (.A(net732),
    .X(net730),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout729 (.A(net732),
    .X(net729),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2259_  (.S0(net1012),
    .A0(\i_ibex/ex_block_i/alu_i/_0110_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0111_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0112_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0113_ ),
    .S1(net1016),
    .X(\i_ibex/ex_block_i/alu_i/_0116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2260_  (.S0(net486),
    .A0(net571),
    .A1(net570),
    .A2(net567),
    .A3(net569),
    .S1(net1208),
    .X(\i_ibex/ex_block_i/alu_i/_0117_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2261_  (.S0(net486),
    .A0(net575),
    .A1(net573),
    .A2(net562),
    .A3(net566),
    .S1(net1208),
    .X(\i_ibex/ex_block_i/alu_i/_0118_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2262_  (.A0(\i_ibex/ex_block_i/alu_i/_0117_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0118_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2263_  (.S0(net486),
    .A0(net579),
    .A1(net577),
    .A2(net556),
    .A3(net559),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0120_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2264_  (.S0(net1050),
    .A0(net554),
    .A1(net552),
    .A2(net591),
    .A3(net594),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2265_  (.A0(\i_ibex/ex_block_i/alu_i/_0120_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0121_ ),
    .S(net1013),
    .X(\i_ibex/ex_block_i/alu_i/_0122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2266_  (.A0(\i_ibex/ex_block_i/alu_i/_0119_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0122_ ),
    .S(net1007),
    .X(\i_ibex/ex_block_i/alu_i/_0123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2267_  (.A(net441),
    .B_N(\i_ibex/ex_block_i/alu_i/_0123_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2268_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net441),
    .A2(\i_ibex/ex_block_i/alu_i/_0116_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0125_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0124_ ));
 sg13g2_buf_2 fanout728 (.A(net732),
    .X(net728),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2270_  (.S0(net1052),
    .A0(net585),
    .A1(net581),
    .A2(net535),
    .A3(net537),
    .S1(net1203),
    .X(\i_ibex/ex_block_i/alu_i/_0127_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2271_  (.S0(net1203),
    .A0(net560),
    .A1(net540),
    .A2(net538),
    .A3(net542),
    .S1(net1052),
    .X(\i_ibex/ex_block_i/alu_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2272_  (.A0(\i_ibex/ex_block_i/alu_i/_0127_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0128_ ),
    .S(net1016),
    .X(\i_ibex/ex_block_i/alu_i/_0129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2273_  (.S0(net486),
    .A0(net546),
    .A1(net544),
    .A2(net531),
    .A3(net534),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2274_  (.S0(net486),
    .A0(net550),
    .A1(net548),
    .A2(net527),
    .A3(net530),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2275_  (.A0(\i_ibex/ex_block_i/alu_i/_0130_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0131_ ),
    .S(net1016),
    .X(\i_ibex/ex_block_i/alu_i/_0132_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2276_  (.A0(\i_ibex/ex_block_i/alu_i/_0129_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0132_ ),
    .S(net1011),
    .X(\i_ibex/ex_block_i/alu_i/_0133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2277_  (.S0(net486),
    .A0(net554),
    .A1(net552),
    .A2(net591),
    .A3(net593),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0134_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2278_  (.S0(net1050),
    .A0(net579),
    .A1(net577),
    .A2(net556),
    .A3(net559),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2279_  (.A0(\i_ibex/ex_block_i/alu_i/_0134_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0135_ ),
    .S(net1013),
    .X(\i_ibex/ex_block_i/alu_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2280_  (.S0(net1050),
    .A0(net575),
    .A1(net573),
    .A2(net562),
    .A3(net565),
    .S1(net1199),
    .X(\i_ibex/ex_block_i/alu_i/_0137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2281_  (.S0(net1050),
    .A0(net571),
    .A1(net570),
    .A2(net567),
    .A3(net569),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0138_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2282_  (.A0(\i_ibex/ex_block_i/alu_i/_0137_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0138_ ),
    .S(net1013),
    .X(\i_ibex/ex_block_i/alu_i/_0139_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2283_  (.A0(\i_ibex/ex_block_i/alu_i/_0136_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0139_ ),
    .S(net1012),
    .X(\i_ibex/ex_block_i/alu_i/_0140_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2284_  (.A0(\i_ibex/ex_block_i/alu_i/_0133_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0140_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2285_  (.A(\i_ibex/ex_block_i/alu_i/_0141_ ),
    .B(net996),
    .Y(\i_ibex/ex_block_i/alu_i/_0142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2286_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0125_ ),
    .A2(net997),
    .Y(\i_ibex/ex_block_i/alu_i/_0143_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0142_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2287_  (.A(net1211),
    .B(\i_ibex/ex_block_i/alu_i/_0143_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2288_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1210),
    .A2(\i_ibex/ex_block_i/alu_i/_0105_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0145_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0144_ ));
 sg13g2_buf_2 fanout727 (.A(net732),
    .X(net727),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout726 (.A(net732),
    .X(net726),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/ex_block_i/alu_i/_2291_  (.B(net1290),
    .A(net1288),
    .X(\i_ibex/ex_block_i/alu_i/_0148_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/ex_block_i/alu_i/_2292_  (.X(\i_ibex/ex_block_i/alu_i/_0149_ ),
    .A(net621),
    .B(\i_ibex/ex_block_i/alu_i/_0064_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0148_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2293_  (.B(\i_ibex/ex_block_i/alu_i/_1290_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0064_ ),
    .A(net1290),
    .Y(\i_ibex/ex_block_i/alu_i/_0150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout725 (.A(net732),
    .X(net725),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 \i_ibex/ex_block_i/alu_i/_2295_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0152_ ),
    .B(net1164),
    .A(net1173));
 sg13g2_buf_2 fanout724 (.A(net732),
    .X(net724),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2297_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net584),
    .A2(net1145),
    .Y(\i_ibex/ex_block_i/alu_i/_0154_ ),
    .B1(\i_ibex/alu_operand_b_ex [31]));
 sg13g2_buf_2 fanout723 (.A(net733),
    .X(net723),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2299_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0156_ ),
    .B(net1169),
    .A(net584));
 sg13g2_buf_2 fanout722 (.A(net733),
    .X(net722),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2301_  (.B(\i_ibex/alu_operand_b_ex [31]),
    .C(net1170),
    .A(net584),
    .Y(\i_ibex/ex_block_i/alu_i/_0158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout721 (.A(\i_ibex/instr_rdata_id [3]),
    .X(net721),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2303_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0156_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0158_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0160_ ),
    .B1(net1175));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2304_  (.A(net1216),
    .B(\i_ibex/ex_block_i/alu_i/_0154_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0160_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2305_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0145_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0161_ ),
    .B1(net1181),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [32]),
    .Y(\i_ibex/ex_block_i/alu_i/_0162_ ),
    .A2(net1150));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2306_  (.A(net1112),
    .B(\i_ibex/ex_block_i/alu_i/_0162_ ),
    .Y(\i_ibex/result_ex [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout720 (.A(net721),
    .X(net720),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/ex_block_i/alu_i/_2308_  (.Y(\i_ibex/ex_block_i/alu_i/_0164_ ),
    .A(net996),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(net721),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout718 (.A(\i_ibex/instr_rdata_id [4]),
    .X(net718),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2312_  (.B(net1011),
    .C(net439),
    .A(net1017),
    .Y(\i_ibex/ex_block_i/alu_i/_0168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2313_  (.A0(\i_ibex/ex_block_i/alu_i/_0127_ ),
    .A1(net1086),
    .S(\i_ibex/ex_block_i/alu_i/_0168_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2314_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0170_ ),
    .B(net1085),
    .A(net996));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2315_  (.B1(\i_ibex/ex_block_i/alu_i/_0170_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0171_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0164_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0169_ ));
 sg13g2_buf_2 fanout716 (.A(net717),
    .X(net716),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout715 (.A(net717),
    .X(net715),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2318_  (.S0(net1050),
    .A0(net552),
    .A1(net550),
    .A2(net593),
    .A3(net528),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0174_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2319_  (.S0(net1051),
    .A0(net544),
    .A1(net542),
    .A2(net533),
    .A3(net539),
    .S1(net1199),
    .X(\i_ibex/ex_block_i/alu_i/_0175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2320_  (.S0(net1051),
    .A0(net548),
    .A1(net546),
    .A2(net529),
    .A3(net532),
    .S1(net1199),
    .X(\i_ibex/ex_block_i/alu_i/_0176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2321_  (.S0(net487),
    .A0(net581),
    .A1(net560),
    .A2(net536),
    .A3(net541),
    .S1(net1209),
    .X(\i_ibex/ex_block_i/alu_i/_0177_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout714 (.A(\i_ibex/instr_rdata_id [5]),
    .X(net714),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2323_  (.S0(net1007),
    .A0(\i_ibex/ex_block_i/alu_i/_0174_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0175_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0176_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0177_ ),
    .S1(net1013),
    .X(\i_ibex/ex_block_i/alu_i/_0179_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout713 (.A(net714),
    .X(net713),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/ex_block_i/alu_i/_2325_  (.Y(\i_ibex/ex_block_i/alu_i/_0181_ ),
    .A(net488),
    .B(net1201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2326_  (.A0(net570),
    .A1(net569),
    .S(\i_ibex/ex_block_i/alu_i/_0181_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0182_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2327_  (.S0(net487),
    .A0(net573),
    .A1(net571),
    .A2(net565),
    .A3(net568),
    .S1(net1208),
    .X(\i_ibex/ex_block_i/alu_i/_0183_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout712 (.A(net714),
    .X(net712),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2329_  (.A0(\i_ibex/ex_block_i/alu_i/_0182_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0183_ ),
    .S(net1018),
    .X(\i_ibex/ex_block_i/alu_i/_0185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2330_  (.S0(net487),
    .A0(net577),
    .A1(net575),
    .A2(net558),
    .A3(net563),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0186_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2331_  (.S0(net1206),
    .A0(net579),
    .A1(net556),
    .A2(net591),
    .A3(net555),
    .S1(net1050),
    .X(\i_ibex/ex_block_i/alu_i/_0187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2332_  (.A0(\i_ibex/ex_block_i/alu_i/_0186_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0187_ ),
    .S(net1018),
    .X(\i_ibex/ex_block_i/alu_i/_0188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2333_  (.A0(\i_ibex/ex_block_i/alu_i/_0185_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0188_ ),
    .S(net1008),
    .X(\i_ibex/ex_block_i/alu_i/_0189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2334_  (.A(net442),
    .B_N(\i_ibex/ex_block_i/alu_i/_0189_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2335_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net442),
    .A2(\i_ibex/ex_block_i/alu_i/_0179_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0191_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0190_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2336_  (.B1(\i_ibex/ex_block_i/alu_i/_0090_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0192_ ),
    .VSS(VSS),
    .A1(net1052),
    .A2(\i_ibex/ex_block_i/alu_i/_0091_ ));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2337_  (.S0(net1052),
    .A0(net581),
    .A1(net560),
    .A2(net536),
    .A3(net540),
    .S1(net1203),
    .X(\i_ibex/ex_block_i/alu_i/_0193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2338_  (.Y(\i_ibex/ex_block_i/alu_i/_0194_ ),
    .A(net1017),
    .B(\i_ibex/ex_block_i/alu_i/_0193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2339_  (.B1(\i_ibex/ex_block_i/alu_i/_0194_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0195_ ),
    .VSS(VSS),
    .A1(net1017),
    .A2(\i_ibex/ex_block_i/alu_i/_0192_ ));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2340_  (.S0(net486),
    .A0(net544),
    .A1(net542),
    .A2(net533),
    .A3(net538),
    .S1(net1209),
    .X(\i_ibex/ex_block_i/alu_i/_0196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2341_  (.S0(net487),
    .A0(net548),
    .A1(net546),
    .A2(net529),
    .A3(net532),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2342_  (.A0(\i_ibex/ex_block_i/alu_i/_0196_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0197_ ),
    .S(net1017),
    .X(\i_ibex/ex_block_i/alu_i/_0198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2343_  (.A0(\i_ibex/ex_block_i/alu_i/_0195_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0198_ ),
    .S(net1011),
    .X(\i_ibex/ex_block_i/alu_i/_0199_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2344_  (.S0(net486),
    .A0(net552),
    .A1(net550),
    .A2(net593),
    .A3(net528),
    .S1(net1206),
    .X(\i_ibex/ex_block_i/alu_i/_0200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2345_  (.S0(net1198),
    .A0(net579),
    .A1(net556),
    .A2(net591),
    .A3(net554),
    .S1(net490),
    .X(\i_ibex/ex_block_i/alu_i/_0201_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2346_  (.A0(\i_ibex/ex_block_i/alu_i/_0200_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0201_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2347_  (.S0(net1050),
    .A0(net577),
    .A1(net575),
    .A2(net558),
    .A3(net563),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2348_  (.S0(net1051),
    .A0(net573),
    .A1(net571),
    .A2(net565),
    .A3(net568),
    .S1(net1198),
    .X(\i_ibex/ex_block_i/alu_i/_0204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2349_  (.A0(\i_ibex/ex_block_i/alu_i/_0203_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0204_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout711 (.A(\i_ibex/instr_rdata_id [6]),
    .X(net711),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2351_  (.A0(\i_ibex/ex_block_i/alu_i/_0202_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0205_ ),
    .S(net1009),
    .X(\i_ibex/ex_block_i/alu_i/_0207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2352_  (.A0(\i_ibex/ex_block_i/alu_i/_0199_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0207_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0208_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2353_  (.A(net994),
    .B(\i_ibex/ex_block_i/alu_i/_0208_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2354_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net994),
    .A2(\i_ibex/ex_block_i/alu_i/_0191_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0210_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0209_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2355_  (.Y(\i_ibex/ex_block_i/alu_i/_0211_ ),
    .A(net1204),
    .B(\i_ibex/ex_block_i/alu_i/_0210_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2356_  (.B1(\i_ibex/ex_block_i/alu_i/_0211_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0212_ ),
    .VSS(VSS),
    .A1(net1204),
    .A2(\i_ibex/ex_block_i/alu_i/_0171_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2357_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net581),
    .A2(net1145),
    .Y(\i_ibex/ex_block_i/alu_i/_0213_ ),
    .B1(\i_ibex/alu_operand_b_ex [30]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2358_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0214_ ),
    .B(net1169),
    .A(net581));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2359_  (.B(\i_ibex/alu_operand_b_ex [30]),
    .C(net1169),
    .A(net581),
    .Y(\i_ibex/ex_block_i/alu_i/_0215_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2360_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0214_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0215_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0216_ ),
    .B1(net1175));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2361_  (.A(net1216),
    .B(\i_ibex/ex_block_i/alu_i/_0213_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0216_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0217_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2362_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0212_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0217_ ),
    .B1(net1180),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [31]),
    .Y(\i_ibex/ex_block_i/alu_i/_0218_ ),
    .A2(net1149));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2363_  (.A(net1112),
    .B(\i_ibex/ex_block_i/alu_i/_0218_ ),
    .Y(\i_ibex/result_ex [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2364_  (.A0(net1085),
    .A1(\i_ibex/ex_block_i/alu_i/_0127_ ),
    .S(net1017),
    .X(\i_ibex/ex_block_i/alu_i/_0219_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2365_  (.A0(\i_ibex/ex_block_i/alu_i/_0128_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0130_ ),
    .S(net1016),
    .X(\i_ibex/ex_block_i/alu_i/_0220_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2366_  (.A0(\i_ibex/ex_block_i/alu_i/_0219_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0220_ ),
    .S(net1011),
    .X(\i_ibex/ex_block_i/alu_i/_0221_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2367_  (.A0(\i_ibex/ex_block_i/alu_i/_0131_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0134_ ),
    .S(net1014),
    .X(\i_ibex/ex_block_i/alu_i/_0222_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2368_  (.A0(\i_ibex/ex_block_i/alu_i/_0135_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0137_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2369_  (.A0(\i_ibex/ex_block_i/alu_i/_0222_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0223_ ),
    .S(net1009),
    .X(\i_ibex/ex_block_i/alu_i/_0224_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2370_  (.A0(\i_ibex/ex_block_i/alu_i/_0138_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0117_ ),
    .S(net1014),
    .X(\i_ibex/ex_block_i/alu_i/_0225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2371_  (.A0(\i_ibex/ex_block_i/alu_i/_0118_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0120_ ),
    .S(net1013),
    .X(\i_ibex/ex_block_i/alu_i/_0226_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2372_  (.A0(\i_ibex/ex_block_i/alu_i/_0225_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0226_ ),
    .S(net1010),
    .X(\i_ibex/ex_block_i/alu_i/_0227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout710 (.A(net711),
    .X(net710),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2374_  (.S0(net440),
    .A0(net1087),
    .A1(\i_ibex/ex_block_i/alu_i/_0221_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0224_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0227_ ),
    .S1(net997),
    .X(\i_ibex/ex_block_i/alu_i/_0229_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2375_  (.A0(net1086),
    .A1(\i_ibex/ex_block_i/alu_i/_0195_ ),
    .S(\i_ibex/ex_block_i/alu_i/_0098_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0230_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2376_  (.A0(\i_ibex/ex_block_i/alu_i/_0198_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0202_ ),
    .S(net1011),
    .X(\i_ibex/ex_block_i/alu_i/_0231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2377_  (.A0(\i_ibex/ex_block_i/alu_i/_0230_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0231_ ),
    .S(net439),
    .X(\i_ibex/ex_block_i/alu_i/_0232_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2378_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0233_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0232_ ),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2379_  (.A(net994),
    .B(net1087),
    .Y(\i_ibex/ex_block_i/alu_i/_0234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2380_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net993),
    .A2(\i_ibex/ex_block_i/alu_i/_0233_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0235_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0234_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2381_  (.A0(\i_ibex/ex_block_i/alu_i/_0229_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0235_ ),
    .S(net1208),
    .X(\i_ibex/ex_block_i/alu_i/_0236_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2382_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net579),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0237_ ),
    .B1(\i_ibex/alu_operand_b_ex [21]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2383_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0238_ ),
    .B(net1168),
    .A(net579));
 sg13g2_buf_2 fanout709 (.A(net710),
    .X(net709),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2385_  (.Y(\i_ibex/ex_block_i/alu_i/_0240_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1046_ ),
    .B(net1168),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2386_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0238_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0240_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0241_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2387_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0237_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0241_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2388_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0236_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0242_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [22]),
    .Y(\i_ibex/ex_block_i/alu_i/_0243_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2389_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0243_ ),
    .Y(\i_ibex/result_ex [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout708 (.A(net710),
    .X(net708),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2391_  (.A0(net1085),
    .A1(\i_ibex/ex_block_i/alu_i/_0129_ ),
    .S(net1011),
    .X(\i_ibex/ex_block_i/alu_i/_0245_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2392_  (.A0(\i_ibex/ex_block_i/alu_i/_0132_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0136_ ),
    .S(net1012),
    .X(\i_ibex/ex_block_i/alu_i/_0246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2393_  (.A0(\i_ibex/ex_block_i/alu_i/_0245_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0246_ ),
    .S(net439),
    .X(\i_ibex/ex_block_i/alu_i/_0247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/ex_block_i/alu_i/_2394_  (.A(\i_ibex/ex_block_i/alu_i/_0164_ ),
    .B(net1085),
    .X(\i_ibex/ex_block_i/alu_i/_0248_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2395_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net995),
    .A2(\i_ibex/ex_block_i/alu_i/_0247_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0249_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ));
 sg13g2_buf_1 fanout707 (.A(\i_ibex/instr_valid_id ),
    .X(net707),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2397_  (.A0(\i_ibex/ex_block_i/alu_i/_0204_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0182_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2398_  (.A0(\i_ibex/ex_block_i/alu_i/_0183_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0186_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0252_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2399_  (.A0(\i_ibex/ex_block_i/alu_i/_0251_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0252_ ),
    .S(net1008),
    .X(\i_ibex/ex_block_i/alu_i/_0253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2400_  (.A0(\i_ibex/ex_block_i/alu_i/_0197_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0200_ ),
    .S(net1014),
    .X(\i_ibex/ex_block_i/alu_i/_0254_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2401_  (.A0(\i_ibex/ex_block_i/alu_i/_0201_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0203_ ),
    .S(net1015),
    .X(\i_ibex/ex_block_i/alu_i/_0255_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2402_  (.A0(\i_ibex/ex_block_i/alu_i/_0254_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0255_ ),
    .S(net1007),
    .X(\i_ibex/ex_block_i/alu_i/_0256_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2403_  (.A(net442),
    .B_N(\i_ibex/ex_block_i/alu_i/_0256_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0257_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2404_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net443),
    .A2(\i_ibex/ex_block_i/alu_i/_0253_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0258_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0257_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2405_  (.B1(\i_ibex/ex_block_i/alu_i/_0090_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0259_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0096_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0091_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2406_  (.A0(\i_ibex/ex_block_i/alu_i/_0193_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0196_ ),
    .S(net1016),
    .X(\i_ibex/ex_block_i/alu_i/_0260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2407_  (.Y(\i_ibex/ex_block_i/alu_i/_0261_ ),
    .A(net1012),
    .B(\i_ibex/ex_block_i/alu_i/_0260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2408_  (.B1(\i_ibex/ex_block_i/alu_i/_0261_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0262_ ),
    .VSS(VSS),
    .A1(net1012),
    .A2(\i_ibex/ex_block_i/alu_i/_0259_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2409_  (.A0(net1087),
    .A1(\i_ibex/ex_block_i/alu_i/_0262_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0263_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2410_  (.A(net992),
    .B(\i_ibex/ex_block_i/alu_i/_0263_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2411_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net992),
    .A2(\i_ibex/ex_block_i/alu_i/_0258_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0265_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0264_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2412_  (.A(net1207),
    .B(\i_ibex/ex_block_i/alu_i/_0265_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2413_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1207),
    .A2(\i_ibex/ex_block_i/alu_i/_0249_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0267_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0266_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2414_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net577),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0268_ ),
    .B1(\i_ibex/alu_operand_b_ex [20]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2415_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0269_ ),
    .B(net1166),
    .A(net577));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2416_  (.Y(\i_ibex/ex_block_i/alu_i/_0270_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1032_ ),
    .B(net1166),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2417_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0269_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0270_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0271_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2418_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0268_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0271_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0272_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2419_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0267_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0272_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [21]),
    .Y(\i_ibex/ex_block_i/alu_i/_0273_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2420_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0273_ ),
    .Y(\i_ibex/result_ex [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2421_  (.A0(\i_ibex/ex_block_i/alu_i/_0139_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0119_ ),
    .S(net1010),
    .X(\i_ibex/ex_block_i/alu_i/_0274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2422_  (.A(net442),
    .B_N(\i_ibex/ex_block_i/alu_i/_0246_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0275_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2423_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net443),
    .A2(\i_ibex/ex_block_i/alu_i/_0274_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0276_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0275_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2424_  (.Y(\i_ibex/ex_block_i/alu_i/_0277_ ),
    .A(net1011),
    .B(net439),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2425_  (.A0(\i_ibex/ex_block_i/alu_i/_0129_ ),
    .A1(net1085),
    .S(\i_ibex/ex_block_i/alu_i/_0277_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2426_  (.A(net996),
    .B(\i_ibex/ex_block_i/alu_i/_0278_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0279_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2427_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net995),
    .A2(\i_ibex/ex_block_i/alu_i/_0276_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0280_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0279_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2428_  (.A0(\i_ibex/ex_block_i/alu_i/_0262_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0256_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0281_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2429_  (.A2(\i_ibex/ex_block_i/alu_i/_0281_ ),
    .A1(net992),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0282_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2430_  (.A0(\i_ibex/ex_block_i/alu_i/_0280_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0282_ ),
    .S(net1207),
    .X(\i_ibex/ex_block_i/alu_i/_0283_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2431_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net575),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0284_ ),
    .B1(\i_ibex/alu_operand_b_ex [19]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2432_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0285_ ),
    .B(net1166),
    .A(net575));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2433_  (.Y(\i_ibex/ex_block_i/alu_i/_0286_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1026_ ),
    .B(net1166),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2434_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0285_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0286_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0287_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2435_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0284_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0287_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0288_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2436_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0283_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0288_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [20]),
    .Y(\i_ibex/ex_block_i/alu_i/_0289_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2437_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0289_ ),
    .Y(\i_ibex/result_ex [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2438_  (.A0(\i_ibex/ex_block_i/alu_i/_0221_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0224_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0290_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2439_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net994),
    .A2(\i_ibex/ex_block_i/alu_i/_0290_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0291_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2440_  (.A0(\i_ibex/ex_block_i/alu_i/_0195_ ),
    .A1(net1085),
    .S(\i_ibex/ex_block_i/alu_i/_0277_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0292_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2441_  (.A0(\i_ibex/ex_block_i/alu_i/_0205_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0185_ ),
    .S(net1008),
    .X(\i_ibex/ex_block_i/alu_i/_0293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2442_  (.A0(\i_ibex/ex_block_i/alu_i/_0231_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0293_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0294_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2443_  (.A0(\i_ibex/ex_block_i/alu_i/_0292_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0294_ ),
    .S(net997),
    .X(\i_ibex/ex_block_i/alu_i/_0295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2444_  (.A(net1211),
    .B(\i_ibex/ex_block_i/alu_i/_0295_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2445_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1210),
    .A2(\i_ibex/ex_block_i/alu_i/_0291_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0297_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0296_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2446_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net573),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0298_ ),
    .B1(\i_ibex/alu_operand_b_ex [18]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2447_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0299_ ),
    .B(net1167),
    .A(net573));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2448_  (.B(\i_ibex/alu_operand_b_ex [18]),
    .C(net1167),
    .A(net573),
    .Y(\i_ibex/ex_block_i/alu_i/_0300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2449_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0299_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0300_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0301_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2450_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0298_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0301_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2451_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0297_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0302_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [19]),
    .Y(\i_ibex/ex_block_i/alu_i/_0303_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2452_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0303_ ),
    .Y(\i_ibex/result_ex [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2453_  (.A0(\i_ibex/ex_block_i/alu_i/_0223_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0225_ ),
    .S(net1009),
    .X(\i_ibex/ex_block_i/alu_i/_0304_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2454_  (.A0(\i_ibex/ex_block_i/alu_i/_0220_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0222_ ),
    .S(net1009),
    .X(\i_ibex/ex_block_i/alu_i/_0305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2455_  (.A(net442),
    .B_N(\i_ibex/ex_block_i/alu_i/_0305_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0306_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2456_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net443),
    .A2(\i_ibex/ex_block_i/alu_i/_0304_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0307_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0306_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2457_  (.A(net996),
    .B(\i_ibex/ex_block_i/alu_i/_0169_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0308_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2458_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net994),
    .A2(\i_ibex/ex_block_i/alu_i/_0307_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0309_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0308_ ));
 sg13g2_inv_1 \i_ibex/ex_block_i/alu_i/_2459_  (.VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0310_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0208_ ),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2460_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net993),
    .A2(\i_ibex/ex_block_i/alu_i/_0310_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0311_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0234_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2461_  (.A0(\i_ibex/ex_block_i/alu_i/_0309_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0311_ ),
    .S(net1210),
    .X(\i_ibex/ex_block_i/alu_i/_0312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2462_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net571),
    .A2(net1145),
    .Y(\i_ibex/ex_block_i/alu_i/_0313_ ),
    .B1(\i_ibex/alu_operand_b_ex [17]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2463_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0314_ ),
    .B(net1169),
    .A(net571));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2464_  (.B(\i_ibex/alu_operand_b_ex [17]),
    .C(net1169),
    .A(net571),
    .Y(\i_ibex/ex_block_i/alu_i/_0315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2465_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0314_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0315_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0316_ ),
    .B1(net1175));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2466_  (.A(net1216),
    .B(\i_ibex/ex_block_i/alu_i/_0313_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0316_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0317_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2467_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0312_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0317_ ),
    .B1(net1180),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [18]),
    .Y(\i_ibex/ex_block_i/alu_i/_0318_ ),
    .A2(net1149));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2468_  (.A(net1112),
    .B(\i_ibex/ex_block_i/alu_i/_0318_ ),
    .Y(\i_ibex/result_ex [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2469_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0141_ ),
    .A2(net997),
    .Y(\i_ibex/ex_block_i/alu_i/_0319_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2470_  (.A0(\i_ibex/ex_block_i/alu_i/_0260_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0254_ ),
    .S(net1012),
    .X(\i_ibex/ex_block_i/alu_i/_0320_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2471_  (.A0(\i_ibex/ex_block_i/alu_i/_0255_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0251_ ),
    .S(net1008),
    .X(\i_ibex/ex_block_i/alu_i/_0321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2472_  (.S0(net440),
    .A0(net1086),
    .A1(\i_ibex/ex_block_i/alu_i/_0102_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0320_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0321_ ),
    .S1(net997),
    .X(\i_ibex/ex_block_i/alu_i/_0322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2473_  (.A(net1210),
    .B(\i_ibex/ex_block_i/alu_i/_0322_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2474_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1210),
    .A2(\i_ibex/ex_block_i/alu_i/_0319_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0324_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0323_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2475_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net570),
    .A2(net1145),
    .Y(\i_ibex/ex_block_i/alu_i/_0325_ ),
    .B1(\i_ibex/alu_operand_b_ex [16]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2476_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0326_ ),
    .B(net1169),
    .A(net570));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2477_  (.B(\i_ibex/alu_operand_b_ex [16]),
    .C(net1169),
    .A(net570),
    .Y(\i_ibex/ex_block_i/alu_i/_0327_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2478_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0326_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0327_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0328_ ),
    .B1(net1175));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2479_  (.A(net1216),
    .B(\i_ibex/ex_block_i/alu_i/_0325_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0328_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2480_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0324_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0329_ ),
    .B1(net1180),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [17]),
    .Y(\i_ibex/ex_block_i/alu_i/_0330_ ),
    .A2(net1149));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2481_  (.A(net1112),
    .B(\i_ibex/ex_block_i/alu_i/_0330_ ),
    .Y(\i_ibex/result_ex [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2482_  (.A(net1204),
    .B(\i_ibex/ex_block_i/alu_i/_0322_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0331_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2483_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1204),
    .A2(\i_ibex/ex_block_i/alu_i/_0319_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0332_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0331_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2484_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net569),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0333_ ),
    .B1(\i_ibex/alu_operand_b_ex [15]));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(net707),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout705 (.A(net706),
    .X(net705),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2487_  (.A(net569),
    .B(net1167),
    .Y(\i_ibex/ex_block_i/alu_i/_0336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2488_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1012_ ),
    .A2(net1167),
    .Y(\i_ibex/ex_block_i/alu_i/_0337_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0336_ ));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2489_  (.B1(\i_ibex/ex_block_i/alu_i/_0071_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0338_ ),
    .VSS(VSS),
    .A1(net1175),
    .A2(\i_ibex/ex_block_i/alu_i/_0337_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2490_  (.A(\i_ibex/ex_block_i/alu_i/_0333_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0338_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0339_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2491_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0332_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0339_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [16]),
    .Y(\i_ibex/ex_block_i/alu_i/_0340_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2492_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0340_ ),
    .Y(\i_ibex/result_ex [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net707),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2494_  (.A0(\i_ibex/ex_block_i/alu_i/_0309_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0311_ ),
    .S(net1205),
    .X(\i_ibex/ex_block_i/alu_i/_0342_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout703 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy [0]),
    .X(net703),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2496_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net567),
    .A2(net1142),
    .Y(\i_ibex/ex_block_i/alu_i/_0344_ ),
    .B1(\i_ibex/alu_operand_b_ex [14]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2497_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0345_ ),
    .B(net1162),
    .A(net567));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2498_  (.B(\i_ibex/alu_operand_b_ex [14]),
    .C(net1163),
    .A(net567),
    .Y(\i_ibex/ex_block_i/alu_i/_0346_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2499_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0345_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0346_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0347_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2500_  (.A(net1213),
    .B(\i_ibex/ex_block_i/alu_i/_0344_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0347_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0348_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2501_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0342_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0348_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [15]),
    .Y(\i_ibex/ex_block_i/alu_i/_0349_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2502_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0349_ ),
    .Y(\i_ibex/result_ex [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout702 (.A(net703),
    .X(net702),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(net703),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(net703),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2506_  (.A(net1205),
    .B(\i_ibex/ex_block_i/alu_i/_0295_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0353_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2507_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1204),
    .A2(\i_ibex/ex_block_i/alu_i/_0291_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0354_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0353_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2508_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net565),
    .A2(net1142),
    .Y(\i_ibex/ex_block_i/alu_i/_0355_ ),
    .B1(\i_ibex/alu_operand_b_ex [13]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2509_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0356_ ),
    .B(net1162),
    .A(net565));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2510_  (.B(\i_ibex/alu_operand_b_ex [13]),
    .C(net1162),
    .A(net565),
    .Y(\i_ibex/ex_block_i/alu_i/_0357_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(net703),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2512_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0356_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0357_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0359_ ),
    .B1(net1172));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2513_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0355_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0359_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0360_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2514_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0354_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0360_ ),
    .B1(net1178),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [14]),
    .Y(\i_ibex/ex_block_i/alu_i/_0361_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2515_  (.A(net1109),
    .B(\i_ibex/ex_block_i/alu_i/_0361_ ),
    .Y(\i_ibex/result_ex [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2516_  (.A0(\i_ibex/ex_block_i/alu_i/_0280_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0282_ ),
    .S(net1200),
    .X(\i_ibex/ex_block_i/alu_i/_0362_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(net703),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2518_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net562),
    .A2(net1142),
    .Y(\i_ibex/ex_block_i/alu_i/_0364_ ),
    .B1(\i_ibex/alu_operand_b_ex [12]));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(\i_ibex/instr_first_cycle_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2520_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0366_ ),
    .B(net1162),
    .A(net562));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2521_  (.B(net1107),
    .C(net1162),
    .A(net562),
    .Y(\i_ibex/ex_block_i/alu_i/_0367_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2522_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0366_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0367_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0368_ ),
    .B1(net1172));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2523_  (.A(net1213),
    .B(\i_ibex/ex_block_i/alu_i/_0364_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0368_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0369_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2524_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0362_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0369_ ),
    .B1(net1178),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [13]),
    .Y(\i_ibex/ex_block_i/alu_i/_0370_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2525_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0370_ ),
    .Y(\i_ibex/result_ex [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2526_  (.S0(net1007),
    .A0(\i_ibex/ex_block_i/alu_i/_0121_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0112_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0110_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0111_ ),
    .S1(net1016),
    .X(\i_ibex/ex_block_i/alu_i/_0371_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2527_  (.A(net441),
    .B_N(\i_ibex/ex_block_i/alu_i/_0227_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2528_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net443),
    .A2(\i_ibex/ex_block_i/alu_i/_0371_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0373_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0372_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2529_  (.A(net997),
    .B(\i_ibex/ex_block_i/alu_i/_0290_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0374_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2530_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net996),
    .A2(\i_ibex/ex_block_i/alu_i/_0373_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0375_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0374_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2531_  (.A2(\i_ibex/ex_block_i/alu_i/_0292_ ),
    .A1(net996),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0376_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2532_  (.A0(\i_ibex/ex_block_i/alu_i/_0375_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0376_ ),
    .S(net1210),
    .X(\i_ibex/ex_block_i/alu_i/_0377_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2533_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net560),
    .A2(net1143),
    .Y(\i_ibex/ex_block_i/alu_i/_0378_ ),
    .B1(\i_ibex/alu_operand_b_ex [29]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2534_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0379_ ),
    .B(net1165),
    .A(net560));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2535_  (.B(\i_ibex/alu_operand_b_ex [29]),
    .C(net1165),
    .A(net560),
    .Y(\i_ibex/ex_block_i/alu_i/_0380_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2536_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0379_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0380_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0381_ ),
    .B1(net1176));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2537_  (.A(net1214),
    .B(\i_ibex/ex_block_i/alu_i/_0378_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0381_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0382_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2538_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0377_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0382_ ),
    .B1(net1178),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [30]),
    .Y(\i_ibex/ex_block_i/alu_i/_0383_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2539_  (.A(net1110),
    .B(\i_ibex/ex_block_i/alu_i/_0383_ ),
    .Y(\i_ibex/result_ex [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2540_  (.A(net1200),
    .B(\i_ibex/ex_block_i/alu_i/_0265_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0384_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2541_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1200),
    .A2(\i_ibex/ex_block_i/alu_i/_0249_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0385_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0384_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2542_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net558),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0386_ ),
    .B1(\i_ibex/alu_operand_b_ex [11]));
 sg13g2_buf_2 fanout696 (.A(net697),
    .X(net696),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2544_  (.A0(net558),
    .A1(\i_ibex/ex_block_i/alu_i/_0908_ ),
    .S(net1162),
    .X(\i_ibex/ex_block_i/alu_i/_0388_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2545_  (.B1(\i_ibex/ex_block_i/alu_i/_0071_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0389_ ),
    .VSS(VSS),
    .A1(net1171),
    .A2(\i_ibex/ex_block_i/alu_i/_0388_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2546_  (.A(\i_ibex/ex_block_i/alu_i/_0386_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0389_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2547_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0385_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0390_ ),
    .B1(net1178),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [12]),
    .Y(\i_ibex/ex_block_i/alu_i/_0391_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2548_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0391_ ),
    .Y(\i_ibex/result_ex [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2549_  (.A0(\i_ibex/ex_block_i/alu_i/_0229_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0235_ ),
    .S(net1201),
    .X(\i_ibex/ex_block_i/alu_i/_0392_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2550_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net556),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0393_ ),
    .B1(\i_ibex/alu_operand_b_ex [10]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2551_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0394_ ),
    .B(net1160),
    .A(net556));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2552_  (.Y(\i_ibex/ex_block_i/alu_i/_0395_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0947_ ),
    .B(net1160),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2553_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0394_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0395_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0396_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2554_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0393_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0396_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2555_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0392_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0397_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [11]),
    .Y(\i_ibex/ex_block_i/alu_i/_0398_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2556_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0398_ ),
    .Y(\i_ibex/result_ex [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2557_  (.A0(\i_ibex/ex_block_i/alu_i/_0127_ ),
    .A1(net1085),
    .S(\i_ibex/ex_block_i/alu_i/_0099_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0399_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2558_  (.A0(\i_ibex/ex_block_i/alu_i/_0399_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0305_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0400_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2559_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net993),
    .A2(\i_ibex/ex_block_i/alu_i/_0400_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0401_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2560_  (.S0(net993),
    .A0(net1087),
    .A1(\i_ibex/ex_block_i/alu_i/_0207_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0199_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0189_ ),
    .S1(net444),
    .X(\i_ibex/ex_block_i/alu_i/_0402_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2561_  (.A(net1200),
    .B(\i_ibex/ex_block_i/alu_i/_0402_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0403_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2562_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1200),
    .A2(\i_ibex/ex_block_i/alu_i/_0401_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0404_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0403_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2563_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net554),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0405_ ),
    .B1(\i_ibex/alu_operand_b_ex [9]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2564_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0406_ ),
    .B(net1162),
    .A(net554));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2565_  (.Y(\i_ibex/ex_block_i/alu_i/_0407_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0938_ ),
    .B(net1162),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2566_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0406_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0407_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0408_ ),
    .B1(net1172));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2567_  (.A(net1213),
    .B(\i_ibex/ex_block_i/alu_i/_0405_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0408_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0409_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2568_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0404_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0409_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [10]),
    .Y(\i_ibex/ex_block_i/alu_i/_0410_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2569_  (.A(net1109),
    .B(\i_ibex/ex_block_i/alu_i/_0410_ ),
    .Y(\i_ibex/result_ex [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2570_  (.A0(\i_ibex/ex_block_i/alu_i/_0102_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0320_ ),
    .S(net438),
    .X(\i_ibex/ex_block_i/alu_i/_0411_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2571_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net994),
    .A2(\i_ibex/ex_block_i/alu_i/_0411_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0412_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2572_  (.S0(\i_ibex/ex_block_i/alu_i/_0164_ ),
    .A0(\i_ibex/ex_block_i/alu_i/_0140_ ),
    .A1(net1085),
    .A2(\i_ibex/ex_block_i/alu_i/_0123_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0133_ ),
    .S1(net444),
    .X(\i_ibex/ex_block_i/alu_i/_0413_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2573_  (.A(net1200),
    .B(\i_ibex/ex_block_i/alu_i/_0413_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0414_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2574_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1200),
    .A2(\i_ibex/ex_block_i/alu_i/_0412_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0415_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0414_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2575_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net552),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0416_ ),
    .B1(\i_ibex/alu_operand_b_ex [8]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2576_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0417_ ),
    .B(net1160),
    .A(net552));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2577_  (.Y(\i_ibex/ex_block_i/alu_i/_0418_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0956_ ),
    .B(net1160),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2578_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0417_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0418_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0419_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2579_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0416_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0419_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0420_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2580_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0415_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0420_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [9]),
    .Y(\i_ibex/ex_block_i/alu_i/_0421_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2581_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0421_ ),
    .Y(\i_ibex/result_ex [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2582_  (.A(net1014),
    .B_N(\i_ibex/ex_block_i/alu_i/_0187_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0422_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2583_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1014),
    .A2(\i_ibex/ex_block_i/alu_i/_0174_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0423_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0422_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2584_  (.A(net1008),
    .B(\i_ibex/ex_block_i/alu_i/_0252_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0424_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2585_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1008),
    .A2(\i_ibex/ex_block_i/alu_i/_0423_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0425_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0424_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2586_  (.A(net441),
    .B_N(\i_ibex/ex_block_i/alu_i/_0321_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0426_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2587_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net443),
    .A2(\i_ibex/ex_block_i/alu_i/_0425_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0427_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0426_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2588_  (.A(net993),
    .B(\i_ibex/ex_block_i/alu_i/_0411_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0428_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2589_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net994),
    .A2(\i_ibex/ex_block_i/alu_i/_0427_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0429_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0428_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2590_  (.A2(\i_ibex/ex_block_i/alu_i/_0088_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0133_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0104_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0430_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/ex_block_i/alu_i/_2591_  (.A0(\i_ibex/ex_block_i/alu_i/_0429_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0430_ ),
    .S(net1201),
    .X(\i_ibex/ex_block_i/alu_i/_0431_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2592_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net550),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0432_ ),
    .B1(\i_ibex/alu_operand_b_ex [7]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2593_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0433_ ),
    .B(net1160),
    .A(net550));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2594_  (.Y(\i_ibex/ex_block_i/alu_i/_0434_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0952_ ),
    .B(net1160),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2595_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0433_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0434_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0435_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2596_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0432_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0435_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0436_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2597_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0431_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0436_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [8]),
    .Y(\i_ibex/ex_block_i/alu_i/_0437_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2598_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0437_ ),
    .Y(\i_ibex/result_ex [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2599_  (.A(net1013),
    .B_N(\i_ibex/ex_block_i/alu_i/_0121_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0438_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2600_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1013),
    .A2(\i_ibex/ex_block_i/alu_i/_0110_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0439_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0438_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2601_  (.A(net1007),
    .B(\i_ibex/ex_block_i/alu_i/_0226_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0440_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2602_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1007),
    .A2(\i_ibex/ex_block_i/alu_i/_0439_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0441_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0440_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2603_  (.A(net441),
    .B_N(\i_ibex/ex_block_i/alu_i/_0304_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0442_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2604_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net443),
    .A2(\i_ibex/ex_block_i/alu_i/_0441_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0443_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0442_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2605_  (.A(net992),
    .B(\i_ibex/ex_block_i/alu_i/_0400_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0444_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2606_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net993),
    .A2(\i_ibex/ex_block_i/alu_i/_0443_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0445_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0444_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2607_  (.A2(\i_ibex/ex_block_i/alu_i/_0199_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0088_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0104_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0446_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2608_  (.A0(\i_ibex/ex_block_i/alu_i/_0445_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0446_ ),
    .S(net1200),
    .X(\i_ibex/ex_block_i/alu_i/_0447_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2609_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net548),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0448_ ),
    .B1(\i_ibex/alu_operand_b_ex [6]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2610_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0449_ ),
    .B(net1160),
    .A(net548));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2611_  (.B(\i_ibex/alu_operand_b_ex [6]),
    .C(net1160),
    .A(net548),
    .Y(\i_ibex/ex_block_i/alu_i/_0450_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2612_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0449_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0450_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0451_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2613_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0448_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0451_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0452_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2614_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0447_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0452_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [7]),
    .Y(\i_ibex/ex_block_i/alu_i/_0453_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2615_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0453_ ),
    .Y(\i_ibex/result_ex [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2616_  (.A(net1014),
    .B_N(\i_ibex/ex_block_i/alu_i/_0174_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0454_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2617_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1014),
    .A2(\i_ibex/ex_block_i/alu_i/_0176_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0455_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0454_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2618_  (.A(net1008),
    .B(\i_ibex/ex_block_i/alu_i/_0188_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0456_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2619_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1008),
    .A2(\i_ibex/ex_block_i/alu_i/_0455_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0457_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0456_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2620_  (.A(net441),
    .B_N(\i_ibex/ex_block_i/alu_i/_0293_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0458_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2621_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net442),
    .A2(\i_ibex/ex_block_i/alu_i/_0457_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0459_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0458_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2622_  (.A(net993),
    .B(\i_ibex/ex_block_i/alu_i/_0232_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0460_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2623_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net993),
    .A2(\i_ibex/ex_block_i/alu_i/_0459_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0461_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0460_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2624_  (.A2(\i_ibex/ex_block_i/alu_i/_0221_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0088_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0104_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0462_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2625_  (.A0(\i_ibex/ex_block_i/alu_i/_0461_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0462_ ),
    .S(net1201),
    .X(\i_ibex/ex_block_i/alu_i/_0463_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2626_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net546),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0464_ ),
    .B1(\i_ibex/alu_operand_b_ex [5]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2627_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0465_ ),
    .B(net1161),
    .A(net546));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2628_  (.Y(\i_ibex/ex_block_i/alu_i/_0466_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0720_ ),
    .B(net1161),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2629_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0465_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0466_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0467_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2630_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0464_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0467_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0468_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2631_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0463_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0468_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [6]),
    .Y(\i_ibex/ex_block_i/alu_i/_0469_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2632_  (.A(net1108),
    .B(\i_ibex/ex_block_i/alu_i/_0469_ ),
    .Y(\i_ibex/result_ex [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout695 (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_110_ ),
    .X(net695),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout694 (.A(\i_ibex/id_stage_i/controller_run ),
    .X(net694),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout693 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0094_ ),
    .X(net693),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2636_  (.A(net1016),
    .B_N(\i_ibex/ex_block_i/alu_i/_0110_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0473_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2637_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1016),
    .A2(\i_ibex/ex_block_i/alu_i/_0112_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0474_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0473_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2638_  (.A(net1007),
    .B(\i_ibex/ex_block_i/alu_i/_0122_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0475_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2639_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1012),
    .A2(\i_ibex/ex_block_i/alu_i/_0474_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0476_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0475_ ));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2640_  (.A(net441),
    .B_N(\i_ibex/ex_block_i/alu_i/_0274_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0477_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2641_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net442),
    .A2(\i_ibex/ex_block_i/alu_i/_0476_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0478_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0477_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2642_  (.A(net995),
    .B(\i_ibex/ex_block_i/alu_i/_0247_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0479_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2643_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net992),
    .A2(\i_ibex/ex_block_i/alu_i/_0478_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0480_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0479_ ));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2644_  (.A2(\i_ibex/ex_block_i/alu_i/_0263_ ),
    .A1(net992),
    .B1(\i_ibex/ex_block_i/alu_i/_0248_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0481_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2645_  (.A0(\i_ibex/ex_block_i/alu_i/_0480_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0481_ ),
    .S(net1203),
    .X(\i_ibex/ex_block_i/alu_i/_0482_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout692 (.A(\i_ibex/csr_op [1]),
    .X(net692),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2647_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net544),
    .A2(net1141),
    .Y(\i_ibex/ex_block_i/alu_i/_0484_ ),
    .B1(\i_ibex/alu_operand_b_ex [4]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2648_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0485_ ),
    .B(net1161),
    .A(net544));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2649_  (.Y(\i_ibex/ex_block_i/alu_i/_0486_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0771_ ),
    .B(net1161),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2650_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0485_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0486_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0487_ ),
    .B1(net1171));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2651_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0484_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0487_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0488_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2652_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0482_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0488_ ),
    .B1(net1177),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [5]),
    .Y(\i_ibex/ex_block_i/alu_i/_0489_ ),
    .A2(net1146));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2653_  (.A(net1109),
    .B(\i_ibex/ex_block_i/alu_i/_0489_ ),
    .Y(\i_ibex/result_ex [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2654_  (.B1(\i_ibex/ex_block_i/alu_i/_0170_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0490_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0164_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0278_ ));
 sg13g2_mux4_1 \i_ibex/ex_block_i/alu_i/_2655_  (.S0(net1007),
    .A0(\i_ibex/ex_block_i/alu_i/_0187_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0176_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0174_ ),
    .A3(\i_ibex/ex_block_i/alu_i/_0175_ ),
    .S1(net1013),
    .X(\i_ibex/ex_block_i/alu_i/_0491_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/ex_block_i/alu_i/_2656_  (.A(net442),
    .B_N(\i_ibex/ex_block_i/alu_i/_0253_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0492_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2657_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net441),
    .A2(\i_ibex/ex_block_i/alu_i/_0491_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0493_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0492_ ));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2658_  (.A(net992),
    .B(\i_ibex/ex_block_i/alu_i/_0281_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0494_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2659_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net992),
    .A2(\i_ibex/ex_block_i/alu_i/_0493_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0495_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0494_ ));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2660_  (.Y(\i_ibex/ex_block_i/alu_i/_0496_ ),
    .A(net1209),
    .B(\i_ibex/ex_block_i/alu_i/_0495_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2661_  (.B1(\i_ibex/ex_block_i/alu_i/_0496_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0497_ ),
    .VSS(VSS),
    .A1(net1209),
    .A2(\i_ibex/ex_block_i/alu_i/_0490_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2662_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net542),
    .A2(\i_ibex/ex_block_i/alu_i/_0152_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0498_ ),
    .B1(\i_ibex/alu_operand_b_ex [3]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2663_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0499_ ),
    .B(net1164),
    .A(net542));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2664_  (.Y(\i_ibex/ex_block_i/alu_i/_0500_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0765_ ),
    .B(net1164),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2665_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0499_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0500_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0501_ ),
    .B1(net1176));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2666_  (.A(net1214),
    .B(\i_ibex/ex_block_i/alu_i/_0498_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0501_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0502_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2667_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0497_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0502_ ),
    .B1(net1181),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [4]),
    .Y(\i_ibex/ex_block_i/alu_i/_0503_ ),
    .A2(net1150));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2668_  (.A(net1110),
    .B(\i_ibex/ex_block_i/alu_i/_0503_ ),
    .Y(\i_ibex/result_ex [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2669_  (.A0(\i_ibex/ex_block_i/alu_i/_0375_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0376_ ),
    .S(net1203),
    .X(\i_ibex/ex_block_i/alu_i/_0504_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2670_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net540),
    .A2(net1143),
    .Y(\i_ibex/ex_block_i/alu_i/_0505_ ),
    .B1(\i_ibex/alu_operand_b_ex [2]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2671_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0506_ ),
    .B(net1164),
    .A(net540));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2672_  (.Y(\i_ibex/ex_block_i/alu_i/_0507_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0780_ ),
    .B(net1164),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2673_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0506_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0507_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0508_ ),
    .B1(net1173));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2674_  (.A(net1214),
    .B(\i_ibex/ex_block_i/alu_i/_0505_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0508_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0509_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2675_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0504_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0509_ ),
    .B1(net1181),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [3]),
    .Y(\i_ibex/ex_block_i/alu_i/_0510_ ),
    .A2(net1150));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2676_  (.A(net1110),
    .B(\i_ibex/ex_block_i/alu_i/_0510_ ),
    .Y(\i_ibex/result_ex [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2677_  (.Y(\i_ibex/ex_block_i/alu_i/_0511_ ),
    .A(net1203),
    .B(\i_ibex/ex_block_i/alu_i/_0495_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2678_  (.B1(\i_ibex/ex_block_i/alu_i/_0511_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0512_ ),
    .VSS(VSS),
    .A1(net1203),
    .A2(\i_ibex/ex_block_i/alu_i/_0490_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2679_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net538),
    .A2(net1143),
    .Y(\i_ibex/ex_block_i/alu_i/_0513_ ),
    .B1(\i_ibex/alu_operand_b_ex [28]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2680_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0514_ ),
    .B(net1165),
    .A(net538));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2681_  (.B(\i_ibex/alu_operand_b_ex [28]),
    .C(net1165),
    .A(net538),
    .Y(\i_ibex/ex_block_i/alu_i/_0515_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2682_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0514_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0515_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0516_ ),
    .B1(net1173));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2683_  (.A(net1214),
    .B(\i_ibex/ex_block_i/alu_i/_0513_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0516_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0517_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2684_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0512_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0517_ ),
    .B1(net1178),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [29]),
    .Y(\i_ibex/ex_block_i/alu_i/_0518_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2685_  (.A(net1110),
    .B(\i_ibex/ex_block_i/alu_i/_0518_ ),
    .Y(\i_ibex/result_ex [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2686_  (.Y(\i_ibex/ex_block_i/alu_i/_0519_ ),
    .A(net1210),
    .B(\i_ibex/ex_block_i/alu_i/_0210_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2687_  (.B1(\i_ibex/ex_block_i/alu_i/_0519_ ),
    .VDD(VDD),
    .Y(\i_ibex/ex_block_i/alu_i/_0520_ ),
    .VSS(VSS),
    .A1(net1209),
    .A2(\i_ibex/ex_block_i/alu_i/_0171_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2688_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net536),
    .A2(net1143),
    .Y(\i_ibex/ex_block_i/alu_i/_0521_ ),
    .B1(net526));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2689_  (.A0(net536),
    .A1(\i_ibex/ex_block_i/alu_i/_0817_ ),
    .S(net1164),
    .X(\i_ibex/ex_block_i/alu_i/_0522_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2690_  (.A(net1173),
    .B(\i_ibex/ex_block_i/alu_i/_0522_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0523_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2691_  (.A(net1213),
    .B(\i_ibex/ex_block_i/alu_i/_0521_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0523_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0524_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2692_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0520_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0524_ ),
    .B1(net1178),
    .A1(net435),
    .Y(\i_ibex/ex_block_i/alu_i/_0525_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2693_  (.A(net1110),
    .B(\i_ibex/ex_block_i/alu_i/_0525_ ),
    .Y(\i_ibex/result_ex [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2694_  (.A0(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .S(net1521),
    .X(\i_ibex/ex_block_i/alu_i/_0526_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/ex_block_i/alu_i/_2695_  (.Y(\i_ibex/ex_block_i/alu_i/_0527_ ),
    .B(\i_ibex/ex_block_i/alu_i/_0526_ ),
    .A_N(net1151),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2696_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1266_ ),
    .A2(net1151),
    .Y(\i_ibex/ex_block_i/alu_i/_0528_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1281_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2697_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1151),
    .A2(\i_ibex/ex_block_i/alu_i/_1300_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0529_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_1295_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2698_  (.A0(\i_ibex/ex_block_i/alu_i/_0528_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0529_ ),
    .S(net1522),
    .X(\i_ibex/ex_block_i/alu_i/_0530_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2699_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_1289_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_1296_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0531_ ),
    .B1(net583));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2700_  (.Y(\i_ibex/ex_block_i/alu_i/_0532_ ),
    .A(\i_ibex/alu_operand_b_ex [31]),
    .B(\i_ibex/ex_block_i/alu_i/_0531_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2701_  (.Y(\i_ibex/ex_block_i/alu_i/_0533_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1304_ ),
    .B(\i_ibex/ex_block_i/alu_i/_1301_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2702_  (.B(\i_ibex/ex_block_i/alu_i/_1299_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0533_ ),
    .A(net583),
    .Y(\i_ibex/ex_block_i/alu_i/_0534_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2703_  (.B(\i_ibex/ex_block_i/alu_i/_0532_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0534_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0611_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0535_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2704_  (.A2(\i_ibex/ex_block_i/alu_i/_0530_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0527_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0535_ ),
    .X(\i_ibex/ex_block_i/alu_i/_0536_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2705_  (.A(net1204),
    .B(\i_ibex/ex_block_i/alu_i/_0143_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0537_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2706_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1204),
    .A2(\i_ibex/ex_block_i/alu_i/_0105_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0538_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0537_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2707_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net535),
    .A2(net1143),
    .Y(\i_ibex/ex_block_i/alu_i/_0539_ ),
    .B1(net488));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2708_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0540_ ),
    .B(net1164),
    .A(net535));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2709_  (.Y(\i_ibex/ex_block_i/alu_i/_0541_ ),
    .A(\i_ibex/ex_block_i/alu_i/_0804_ ),
    .B(net1164),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2710_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0540_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0541_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0542_ ),
    .B1(net1173));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2711_  (.A(net1213),
    .B(\i_ibex/ex_block_i/alu_i/_0539_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0542_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0543_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2712_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0538_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0543_ ),
    .B1(net1180),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [1]),
    .Y(\i_ibex/ex_block_i/alu_i/_0544_ ),
    .A2(net1149));
 sg13g2_a21o_1 \i_ibex/ex_block_i/alu_i/_2713_  (.A2(\i_ibex/ex_block_i/alu_i/_0544_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0536_ ),
    .B1(net1112),
    .X(\i_ibex/ex_block_i/alu_i/_0545_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/ex_block_i/alu_i/_2714_  (.B1(\i_ibex/ex_block_i/alu_i/_0545_ ),
    .VDD(VDD),
    .Y(\i_ibex/result_ex [0]),
    .VSS(VSS),
    .A1(\i_ibex/ex_block_i/alu_i/_0668_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0061_ ));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2715_  (.A0(\i_ibex/ex_block_i/alu_i/_0480_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0481_ ),
    .S(net1209),
    .X(\i_ibex/ex_block_i/alu_i/_0546_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2716_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net533),
    .A2(net1143),
    .Y(\i_ibex/ex_block_i/alu_i/_0547_ ),
    .B1(\i_ibex/alu_operand_b_ex [27]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2717_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0548_ ),
    .B(net1165),
    .A(net533));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2718_  (.B(\i_ibex/alu_operand_b_ex [27]),
    .C(net1165),
    .A(net533),
    .Y(\i_ibex/ex_block_i/alu_i/_0549_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2719_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0548_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0549_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0550_ ),
    .B1(net1173));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2720_  (.A(net1213),
    .B(\i_ibex/ex_block_i/alu_i/_0547_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0550_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0551_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2721_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0546_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0551_ ),
    .B1(net1178),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [28]),
    .Y(\i_ibex/ex_block_i/alu_i/_0552_ ),
    .A2(net1147));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2722_  (.A(net1109),
    .B(\i_ibex/ex_block_i/alu_i/_0552_ ),
    .Y(\i_ibex/result_ex [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2723_  (.A0(\i_ibex/ex_block_i/alu_i/_0461_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0462_ ),
    .S(net1208),
    .X(\i_ibex/ex_block_i/alu_i/_0553_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2724_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net531),
    .A2(net1142),
    .Y(\i_ibex/ex_block_i/alu_i/_0554_ ),
    .B1(\i_ibex/alu_operand_b_ex [26]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2725_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0555_ ),
    .B(net1163),
    .A(net531));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2726_  (.B(\i_ibex/alu_operand_b_ex [26]),
    .C(net1163),
    .A(net531),
    .Y(\i_ibex/ex_block_i/alu_i/_0556_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2727_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0555_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0556_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0557_ ),
    .B1(net1172));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2728_  (.A(net1212),
    .B(\i_ibex/ex_block_i/alu_i/_0554_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0557_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0558_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2729_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0553_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0558_ ),
    .B1(net1180),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [27]),
    .Y(\i_ibex/ex_block_i/alu_i/_0559_ ),
    .A2(net1149));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2730_  (.A(net1112),
    .B(\i_ibex/ex_block_i/alu_i/_0559_ ),
    .Y(\i_ibex/result_ex [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2731_  (.A0(\i_ibex/ex_block_i/alu_i/_0445_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0446_ ),
    .S(net1207),
    .X(\i_ibex/ex_block_i/alu_i/_0560_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2732_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net529),
    .A2(net1145),
    .Y(\i_ibex/ex_block_i/alu_i/_0561_ ),
    .B1(\i_ibex/alu_operand_b_ex [25]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2733_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0562_ ),
    .B(net1166),
    .A(net529));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2734_  (.Y(\i_ibex/ex_block_i/alu_i/_0563_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1065_ ),
    .B(net1166),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2735_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0562_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0563_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0564_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2736_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0561_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0564_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0565_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2737_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0560_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0565_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [26]),
    .Y(\i_ibex/ex_block_i/alu_i/_0566_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2738_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0566_ ),
    .Y(\i_ibex/result_ex [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/ex_block_i/alu_i/_2739_  (.A0(\i_ibex/ex_block_i/alu_i/_0429_ ),
    .A1(\i_ibex/ex_block_i/alu_i/_0430_ ),
    .S(net1208),
    .X(\i_ibex/ex_block_i/alu_i/_0567_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2740_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net527),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0568_ ),
    .B1(\i_ibex/alu_operand_b_ex [24]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2741_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0569_ ),
    .B(net1166),
    .A(net527));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2742_  (.Y(\i_ibex/ex_block_i/alu_i/_0570_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1082_ ),
    .B(net1166),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2743_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0569_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0570_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0571_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2744_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0568_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0571_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0572_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2745_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0567_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0572_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [25]),
    .Y(\i_ibex/ex_block_i/alu_i/_0573_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2746_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0573_ ),
    .Y(\i_ibex/result_ex [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2747_  (.A(net1207),
    .B(\i_ibex/ex_block_i/alu_i/_0413_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0574_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2748_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1207),
    .A2(\i_ibex/ex_block_i/alu_i/_0412_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0575_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0574_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2749_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net593),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0576_ ),
    .B1(\i_ibex/alu_operand_b_ex [23]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2750_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0577_ ),
    .B(net1168),
    .A(net593));
 sg13g2_nand2_1 \i_ibex/ex_block_i/alu_i/_2751_  (.Y(\i_ibex/ex_block_i/alu_i/_0578_ ),
    .A(\i_ibex/ex_block_i/alu_i/_1078_ ),
    .B(net1168),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2752_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0577_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0578_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0579_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2753_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0576_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0579_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0580_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2754_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0575_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0580_ ),
    .B1(net1180),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [24]),
    .Y(\i_ibex/ex_block_i/alu_i/_0581_ ),
    .A2(net1149));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2755_  (.A(net1112),
    .B(\i_ibex/ex_block_i/alu_i/_0581_ ),
    .Y(\i_ibex/result_ex [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2756_  (.A(net1207),
    .B(\i_ibex/ex_block_i/alu_i/_0402_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0582_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2757_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1207),
    .A2(\i_ibex/ex_block_i/alu_i/_0401_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0583_ ),
    .B1(\i_ibex/ex_block_i/alu_i/_0582_ ));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2758_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net592),
    .A2(net1144),
    .Y(\i_ibex/ex_block_i/alu_i/_0584_ ),
    .B1(\i_ibex/alu_operand_b_ex [22]));
 sg13g2_or2_1 \i_ibex/ex_block_i/alu_i/_2759_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/ex_block_i/alu_i/_0585_ ),
    .B(net1168),
    .A(net591));
 sg13g2_nand3_1 \i_ibex/ex_block_i/alu_i/_2760_  (.B(\i_ibex/alu_operand_b_ex [22]),
    .C(net1168),
    .A(net592),
    .Y(\i_ibex/ex_block_i/alu_i/_0586_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/ex_block_i/alu_i/_2761_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_i/_0585_ ),
    .A2(\i_ibex/ex_block_i/alu_i/_0586_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0587_ ),
    .B1(net1174));
 sg13g2_nor3_1 \i_ibex/ex_block_i/alu_i/_2762_  (.A(net1215),
    .B(\i_ibex/ex_block_i/alu_i/_0584_ ),
    .C(\i_ibex/ex_block_i/alu_i/_0587_ ),
    .Y(\i_ibex/ex_block_i/alu_i/_0588_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/ex_block_i/alu_i/_2763_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/ex_block_i/alu_i/_0583_ ),
    .C1(\i_ibex/ex_block_i/alu_i/_0588_ ),
    .B1(net1179),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [23]),
    .Y(\i_ibex/ex_block_i/alu_i/_0589_ ),
    .A2(net1148));
 sg13g2_nor2_1 \i_ibex/ex_block_i/alu_i/_2764_  (.A(net1111),
    .B(\i_ibex/ex_block_i/alu_i/_0589_ ),
    .Y(\i_ibex/result_ex [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1360__322  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net322));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout690 (.A(net692),
    .X(net690),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout689 (.A(net692),
    .X(net689),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_0631_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0359_ ),
    .A(net688),
    .VSS(VSS));
 sg13g2_buf_2 fanout688 (.A(\i_ibex/lsu_addr_incr_req ),
    .X(net688),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_0633_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0361_ ),
    .A(net1299),
    .VSS(VSS));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net688),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0635_  (.X(\i_ibex/id_stage_i/_0363_ ),
    .A(net1380),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0636_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [31]),
    .Y(\i_ibex/id_stage_i/_0364_ ),
    .B1(\i_ibex/id_stage_i/_0363_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0637_  (.Y(\i_ibex/id_stage_i/_0365_ ),
    .A(\i_ibex/id_stage_i/alu_op_a_mux_sel_dec [1]),
    .B(net1377),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/_0638_  (.A(net1296),
    .B(\i_ibex/id_stage_i/_0365_ ),
    .Y(\i_ibex/id_stage_i/_0366_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(net687),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/_0640_  (.A(net1259),
    .B(\i_ibex/id_stage_i/imm_a_mux_sel ),
    .C(\i_ibex/id_stage_i/_0365_ ),
    .Y(\i_ibex/id_stage_i/_0368_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(net687),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(net687),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net687),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0644_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [31]),
    .X(\i_ibex/id_stage_i/_0372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0645_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net328),
    .C1(\i_ibex/id_stage_i/_0372_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [31]),
    .Y(\i_ibex/id_stage_i/_0373_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0646_  (.B1(\i_ibex/id_stage_i/_0373_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [31]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0364_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0647_  (.X(\i_ibex/id_stage_i/_0374_ ),
    .A(net1377),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0648_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1298),
    .A2(\i_ibex/lsu_addr_last [30]),
    .Y(\i_ibex/id_stage_i/_0375_ ),
    .B1(\i_ibex/id_stage_i/_0374_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0649_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [30]),
    .X(\i_ibex/id_stage_i/_0376_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0650_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net329),
    .C1(\i_ibex/id_stage_i/_0376_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [30]),
    .Y(\i_ibex/id_stage_i/_0377_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0651_  (.B1(\i_ibex/id_stage_i/_0377_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [30]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0375_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0652_  (.X(\i_ibex/id_stage_i/_0378_ ),
    .A(net1377),
    .B(net1260),
    .C(\i_ibex/rf_rdata_a [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0653_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [21]),
    .Y(\i_ibex/id_stage_i/_0379_ ),
    .B1(\i_ibex/id_stage_i/_0378_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0654_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [21]),
    .X(\i_ibex/id_stage_i/_0380_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0655_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net330),
    .C1(\i_ibex/id_stage_i/_0380_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [21]),
    .Y(\i_ibex/id_stage_i/_0381_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0656_  (.B1(\i_ibex/id_stage_i/_0381_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [21]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0379_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0657_  (.X(\i_ibex/id_stage_i/_0382_ ),
    .A(net1379),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0658_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1298),
    .A2(\i_ibex/lsu_addr_last [20]),
    .Y(\i_ibex/id_stage_i/_0383_ ),
    .B1(\i_ibex/id_stage_i/_0382_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0659_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [20]),
    .X(\i_ibex/id_stage_i/_0384_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0660_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net331),
    .C1(\i_ibex/id_stage_i/_0384_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [20]),
    .Y(\i_ibex/id_stage_i/_0385_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0661_  (.B1(\i_ibex/id_stage_i/_0385_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [20]),
    .VSS(VSS),
    .A1(net1304),
    .A2(\i_ibex/id_stage_i/_0383_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0662_  (.X(\i_ibex/id_stage_i/_0386_ ),
    .A(net1379),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0663_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [19]),
    .Y(\i_ibex/id_stage_i/_0387_ ),
    .B1(\i_ibex/id_stage_i/_0386_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0664_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [19]),
    .X(\i_ibex/id_stage_i/_0388_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0665_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net332),
    .C1(\i_ibex/id_stage_i/_0388_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [19]),
    .Y(\i_ibex/id_stage_i/_0389_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0666_  (.B1(\i_ibex/id_stage_i/_0389_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [19]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0387_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0667_  (.X(\i_ibex/id_stage_i/_0390_ ),
    .A(net1379),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0668_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [18]),
    .Y(\i_ibex/id_stage_i/_0391_ ),
    .B1(\i_ibex/id_stage_i/_0390_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0669_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [18]),
    .X(\i_ibex/id_stage_i/_0392_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0670_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net333),
    .C1(\i_ibex/id_stage_i/_0392_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [18]),
    .Y(\i_ibex/id_stage_i/_0393_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0671_  (.B1(\i_ibex/id_stage_i/_0393_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [18]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0391_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0672_  (.X(\i_ibex/id_stage_i/_0394_ ),
    .A(net1377),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0673_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1298),
    .A2(\i_ibex/lsu_addr_last [17]),
    .Y(\i_ibex/id_stage_i/_0395_ ),
    .B1(\i_ibex/id_stage_i/_0394_ ));
 sg13g2_buf_2 fanout682 (.A(net687),
    .X(net682),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0675_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [17]),
    .X(\i_ibex/id_stage_i/_0397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0676_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net334),
    .C1(\i_ibex/id_stage_i/_0397_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [17]),
    .Y(\i_ibex/id_stage_i/_0398_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0677_  (.B1(\i_ibex/id_stage_i/_0398_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [17]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0395_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0678_  (.X(\i_ibex/id_stage_i/_0399_ ),
    .A(net1378),
    .B(net1260),
    .C(\i_ibex/rf_rdata_a [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0679_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [16]),
    .Y(\i_ibex/id_stage_i/_0400_ ),
    .B1(\i_ibex/id_stage_i/_0399_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0680_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [16]),
    .X(\i_ibex/id_stage_i/_0401_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0681_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net335),
    .C1(\i_ibex/id_stage_i/_0401_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [16]),
    .Y(\i_ibex/id_stage_i/_0402_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0682_  (.B1(\i_ibex/id_stage_i/_0402_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [16]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0400_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0683_  (.X(\i_ibex/id_stage_i/_0403_ ),
    .A(net1379),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0684_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1298),
    .A2(\i_ibex/lsu_addr_last [15]),
    .Y(\i_ibex/id_stage_i/_0404_ ),
    .B1(\i_ibex/id_stage_i/_0403_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0685_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [15]),
    .X(\i_ibex/id_stage_i/_0405_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0686_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net336),
    .C1(\i_ibex/id_stage_i/_0405_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [15]),
    .Y(\i_ibex/id_stage_i/_0406_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0687_  (.B1(\i_ibex/id_stage_i/_0406_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [15]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0404_ ));
 sg13g2_buf_2 fanout681 (.A(net687),
    .X(net681),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0689_  (.X(\i_ibex/id_stage_i/_0408_ ),
    .A(net1377),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0690_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [14]),
    .Y(\i_ibex/id_stage_i/_0409_ ),
    .B1(\i_ibex/id_stage_i/_0408_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0691_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [14]),
    .X(\i_ibex/id_stage_i/_0410_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0692_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net337),
    .C1(\i_ibex/id_stage_i/_0410_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [14]),
    .Y(\i_ibex/id_stage_i/_0411_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0693_  (.B1(\i_ibex/id_stage_i/_0411_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [14]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0409_ ));
 sg13g2_buf_2 fanout680 (.A(net687),
    .X(net680),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net687),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout678 (.A(\i_ibex/id_stage_i/imm_b_mux_sel_dec [1]),
    .X(net678),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0697_  (.X(\i_ibex/id_stage_i/_0415_ ),
    .A(net1379),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0698_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/_0415_ ),
    .Y(\i_ibex/id_stage_i/_0416_ ),
    .A2(\i_ibex/lsu_addr_last [13]),
    .A1(net1298));
 sg13g2_buf_1 fanout677 (.A(net678),
    .X(net677),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net678),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0701_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [13]),
    .X(\i_ibex/id_stage_i/_0419_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0702_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net338),
    .C1(\i_ibex/id_stage_i/_0419_ ),
    .B1(net1194),
    .A1(\i_ibex/pc_id [13]),
    .Y(\i_ibex/id_stage_i/_0420_ ),
    .A2(net1255));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0703_  (.B1(\i_ibex/id_stage_i/_0420_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [13]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0416_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0704_  (.X(\i_ibex/id_stage_i/_0421_ ),
    .A(net1378),
    .B(net1260),
    .C(\i_ibex/rf_rdata_a [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0705_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1295),
    .A2(\i_ibex/lsu_addr_last [12]),
    .Y(\i_ibex/id_stage_i/_0422_ ),
    .B1(\i_ibex/id_stage_i/_0421_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0706_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [12]),
    .X(\i_ibex/id_stage_i/_0423_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0707_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net339),
    .C1(\i_ibex/id_stage_i/_0423_ ),
    .B1(net1194),
    .A1(\i_ibex/pc_id [12]),
    .Y(\i_ibex/id_stage_i/_0424_ ),
    .A2(net1255));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0708_  (.B1(\i_ibex/id_stage_i/_0424_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [12]),
    .VSS(VSS),
    .A1(net1301),
    .A2(\i_ibex/id_stage_i/_0422_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0709_  (.X(\i_ibex/id_stage_i/_0425_ ),
    .A(net1377),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0710_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1295),
    .A2(\i_ibex/lsu_addr_last [29]),
    .Y(\i_ibex/id_stage_i/_0426_ ),
    .B1(\i_ibex/id_stage_i/_0425_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0711_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [29]),
    .X(\i_ibex/id_stage_i/_0427_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0712_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net340),
    .C1(\i_ibex/id_stage_i/_0427_ ),
    .B1(net1194),
    .A1(\i_ibex/pc_id [29]),
    .Y(\i_ibex/id_stage_i/_0428_ ),
    .A2(net1255));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0713_  (.B1(\i_ibex/id_stage_i/_0428_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [29]),
    .VSS(VSS),
    .A1(net1301),
    .A2(\i_ibex/id_stage_i/_0426_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0714_  (.X(\i_ibex/id_stage_i/_0429_ ),
    .A(net1379),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0715_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1295),
    .A2(\i_ibex/lsu_addr_last [11]),
    .Y(\i_ibex/id_stage_i/_0430_ ),
    .B1(\i_ibex/id_stage_i/_0429_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0716_  (.A(net681),
    .B(\i_ibex/lsu_addr_last [11]),
    .X(\i_ibex/id_stage_i/_0431_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0717_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net341),
    .C1(\i_ibex/id_stage_i/_0431_ ),
    .B1(net1194),
    .A1(\i_ibex/pc_id [11]),
    .Y(\i_ibex/id_stage_i/_0432_ ),
    .A2(net1255));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0718_  (.B1(\i_ibex/id_stage_i/_0432_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [11]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0430_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0719_  (.X(\i_ibex/id_stage_i/_0433_ ),
    .A(net1379),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0720_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [10]),
    .Y(\i_ibex/id_stage_i/_0434_ ),
    .B1(\i_ibex/id_stage_i/_0433_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0721_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [10]),
    .X(\i_ibex/id_stage_i/_0435_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0722_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net342),
    .C1(\i_ibex/id_stage_i/_0435_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [10]),
    .Y(\i_ibex/id_stage_i/_0436_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0723_  (.B1(\i_ibex/id_stage_i/_0436_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [10]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0434_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0724_  (.X(\i_ibex/id_stage_i/_0437_ ),
    .A(net1378),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0725_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1295),
    .A2(\i_ibex/lsu_addr_last [9]),
    .Y(\i_ibex/id_stage_i/_0438_ ),
    .B1(\i_ibex/id_stage_i/_0437_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0726_  (.A(net680),
    .B(\i_ibex/lsu_addr_last [9]),
    .X(\i_ibex/id_stage_i/_0439_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0727_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net343),
    .C1(\i_ibex/id_stage_i/_0439_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [9]),
    .Y(\i_ibex/id_stage_i/_0440_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0728_  (.B1(\i_ibex/id_stage_i/_0440_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [9]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0438_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0729_  (.X(\i_ibex/id_stage_i/_0441_ ),
    .A(net1378),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0730_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [8]),
    .Y(\i_ibex/id_stage_i/_0442_ ),
    .B1(\i_ibex/id_stage_i/_0441_ ));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(net678),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0732_  (.A(net683),
    .B(\i_ibex/lsu_addr_last [8]),
    .X(\i_ibex/id_stage_i/_0444_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0733_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net344),
    .C1(\i_ibex/id_stage_i/_0444_ ),
    .B1(net1195),
    .A1(\i_ibex/pc_id [8]),
    .Y(\i_ibex/id_stage_i/_0445_ ),
    .A2(net1256));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0734_  (.B1(\i_ibex/id_stage_i/_0445_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [8]),
    .VSS(VSS),
    .A1(net1301),
    .A2(\i_ibex/id_stage_i/_0442_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0735_  (.X(\i_ibex/id_stage_i/_0446_ ),
    .A(net1380),
    .B(net1262),
    .C(\i_ibex/rf_rdata_a [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0736_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/_0446_ ),
    .Y(\i_ibex/id_stage_i/_0447_ ),
    .A2(\i_ibex/lsu_addr_last [7]),
    .A1(net1294));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0737_  (.A(net683),
    .B(\i_ibex/lsu_addr_last [7]),
    .X(\i_ibex/id_stage_i/_0448_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0738_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net345),
    .C1(\i_ibex/id_stage_i/_0448_ ),
    .B1(net1195),
    .A1(\i_ibex/pc_id [7]),
    .Y(\i_ibex/id_stage_i/_0449_ ),
    .A2(net1256));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0739_  (.B1(\i_ibex/id_stage_i/_0449_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [7]),
    .VSS(VSS),
    .A1(net1301),
    .A2(\i_ibex/id_stage_i/_0447_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0740_  (.X(\i_ibex/id_stage_i/_0450_ ),
    .A(net1377),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0741_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [6]),
    .Y(\i_ibex/id_stage_i/_0451_ ),
    .B1(\i_ibex/id_stage_i/_0450_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0742_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [6]),
    .X(\i_ibex/id_stage_i/_0452_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0743_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net346),
    .C1(\i_ibex/id_stage_i/_0452_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [6]),
    .Y(\i_ibex/id_stage_i/_0453_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0744_  (.B1(\i_ibex/id_stage_i/_0453_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [6]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0451_ ));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net678),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0746_  (.X(\i_ibex/id_stage_i/_0455_ ),
    .A(net1380),
    .B(net1262),
    .C(\i_ibex/rf_rdata_a [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0747_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [5]),
    .Y(\i_ibex/id_stage_i/_0456_ ),
    .B1(\i_ibex/id_stage_i/_0455_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0748_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [5]),
    .X(\i_ibex/id_stage_i/_0457_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0749_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net347),
    .C1(\i_ibex/id_stage_i/_0457_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [5]),
    .Y(\i_ibex/id_stage_i/_0458_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0750_  (.B1(\i_ibex/id_stage_i/_0458_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [5]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0456_ ));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net678),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout672 (.A(\i_ibex/if_stage_i/fetch_rdata [15]),
    .X(net672),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0754_  (.X(\i_ibex/id_stage_i/_0462_ ),
    .A(\i_ibex/id_stage_i/_0359_ ),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0755_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [4]),
    .Y(\i_ibex/id_stage_i/_0463_ ),
    .B1(\i_ibex/id_stage_i/_0462_ ));
 sg13g2_buf_2 fanout670 (.A(net672),
    .X(net670),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout669 (.A(net672),
    .X(net669),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0758_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [4]),
    .X(\i_ibex/id_stage_i/_0466_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0759_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .C1(\i_ibex/id_stage_i/_0466_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [4]),
    .Y(\i_ibex/id_stage_i/_0467_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0760_  (.B1(\i_ibex/id_stage_i/_0467_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [4]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0463_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0761_  (.X(\i_ibex/id_stage_i/_0468_ ),
    .A(net1380),
    .B(net1262),
    .C(\i_ibex/rf_rdata_a [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0762_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1294),
    .A2(\i_ibex/lsu_addr_last [3]),
    .Y(\i_ibex/id_stage_i/_0469_ ),
    .B1(\i_ibex/id_stage_i/_0468_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0763_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [3]),
    .X(\i_ibex/id_stage_i/_0470_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0764_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .C1(\i_ibex/id_stage_i/_0470_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [3]),
    .Y(\i_ibex/id_stage_i/_0471_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0765_  (.B1(\i_ibex/id_stage_i/_0471_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [3]),
    .VSS(VSS),
    .A1(net1300),
    .A2(\i_ibex/id_stage_i/_0469_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0766_  (.X(\i_ibex/id_stage_i/_0472_ ),
    .A(net1378),
    .B(net1263),
    .C(\i_ibex/rf_rdata_a [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0767_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1296),
    .A2(\i_ibex/lsu_addr_last [2]),
    .Y(\i_ibex/id_stage_i/_0473_ ),
    .B1(\i_ibex/id_stage_i/_0472_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0768_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [2]),
    .X(\i_ibex/id_stage_i/_0474_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0769_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .C1(\i_ibex/id_stage_i/_0474_ ),
    .B1(net1195),
    .A1(\i_ibex/pc_id [2]),
    .Y(\i_ibex/id_stage_i/_0475_ ),
    .A2(net1256));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0770_  (.B1(\i_ibex/id_stage_i/_0475_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [2]),
    .VSS(VSS),
    .A1(net1301),
    .A2(\i_ibex/id_stage_i/_0473_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0771_  (.X(\i_ibex/id_stage_i/_0476_ ),
    .A(net1380),
    .B(net1262),
    .C(\i_ibex/rf_rdata_a [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0772_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1298),
    .A2(\i_ibex/lsu_addr_last [28]),
    .Y(\i_ibex/id_stage_i/_0477_ ),
    .B1(\i_ibex/id_stage_i/_0476_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0773_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [28]),
    .X(\i_ibex/id_stage_i/_0478_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0774_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net348),
    .C1(\i_ibex/id_stage_i/_0478_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [28]),
    .Y(\i_ibex/id_stage_i/_0479_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0775_  (.B1(\i_ibex/id_stage_i/_0479_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [28]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0477_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0776_  (.X(\i_ibex/id_stage_i/_0480_ ),
    .A(net1381),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0777_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/_0480_ ),
    .Y(\i_ibex/id_stage_i/_0481_ ),
    .A2(\i_ibex/lsu_addr_last [1]),
    .A1(net1299));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0778_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [1]),
    .X(\i_ibex/id_stage_i/_0482_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0779_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net766),
    .C1(\i_ibex/id_stage_i/_0482_ ),
    .B1(net1193),
    .A1(\i_ibex/pc_id [1]),
    .Y(\i_ibex/id_stage_i/_0483_ ),
    .A2(net1254));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0780_  (.B1(\i_ibex/id_stage_i/_0483_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [1]),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/alu_op_a_mux_sel_dec [1]),
    .A2(\i_ibex/id_stage_i/_0481_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0781_  (.X(\i_ibex/id_stage_i/_0484_ ),
    .A(net1379),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0782_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/_0484_ ),
    .Y(\i_ibex/id_stage_i/_0485_ ),
    .A2(\i_ibex/lsu_addr_last [0]),
    .A1(net1299));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0783_  (.A(net682),
    .B(\i_ibex/lsu_addr_last [0]),
    .X(\i_ibex/id_stage_i/_0486_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0784_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net768),
    .C1(\i_ibex/id_stage_i/_0486_ ),
    .B1(net1195),
    .A1(\i_ibex/pc_id [0]),
    .Y(\i_ibex/id_stage_i/_0487_ ),
    .A2(net1256));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0785_  (.B1(\i_ibex/id_stage_i/_0487_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [0]),
    .VSS(VSS),
    .A1(net1301),
    .A2(\i_ibex/id_stage_i/_0485_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0786_  (.X(\i_ibex/id_stage_i/_0488_ ),
    .A(net1380),
    .B(net1262),
    .C(\i_ibex/rf_rdata_a [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0787_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1295),
    .A2(\i_ibex/lsu_addr_last [27]),
    .Y(\i_ibex/id_stage_i/_0489_ ),
    .B1(\i_ibex/id_stage_i/_0488_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0788_  (.A(net679),
    .B(\i_ibex/lsu_addr_last [27]),
    .X(\i_ibex/id_stage_i/_0490_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0789_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net349),
    .C1(\i_ibex/id_stage_i/_0490_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [27]),
    .Y(\i_ibex/id_stage_i/_0491_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0790_  (.B1(\i_ibex/id_stage_i/_0491_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [27]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0489_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0791_  (.X(\i_ibex/id_stage_i/_0492_ ),
    .A(net1377),
    .B(net1260),
    .C(\i_ibex/rf_rdata_a [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0792_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [26]),
    .Y(\i_ibex/id_stage_i/_0493_ ),
    .B1(\i_ibex/id_stage_i/_0492_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0793_  (.A(net679),
    .B(\i_ibex/lsu_addr_last [26]),
    .X(\i_ibex/id_stage_i/_0494_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0794_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net350),
    .C1(\i_ibex/id_stage_i/_0494_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [26]),
    .Y(\i_ibex/id_stage_i/_0495_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0795_  (.B1(\i_ibex/id_stage_i/_0495_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [26]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0493_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0796_  (.X(\i_ibex/id_stage_i/_0496_ ),
    .A(net1378),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0797_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1298),
    .A2(\i_ibex/lsu_addr_last [25]),
    .Y(\i_ibex/id_stage_i/_0497_ ),
    .B1(\i_ibex/id_stage_i/_0496_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0798_  (.A(net679),
    .B(\i_ibex/lsu_addr_last [25]),
    .X(\i_ibex/id_stage_i/_0498_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0799_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net351),
    .C1(\i_ibex/id_stage_i/_0498_ ),
    .B1(net1197),
    .A1(\i_ibex/pc_id [25]),
    .Y(\i_ibex/id_stage_i/_0499_ ),
    .A2(net1258));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0800_  (.B1(\i_ibex/id_stage_i/_0499_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [25]),
    .VSS(VSS),
    .A1(net1303),
    .A2(\i_ibex/id_stage_i/_0497_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0801_  (.X(\i_ibex/id_stage_i/_0500_ ),
    .A(net1380),
    .B(net1262),
    .C(\i_ibex/rf_rdata_a [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0802_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [24]),
    .Y(\i_ibex/id_stage_i/_0501_ ),
    .B1(\i_ibex/id_stage_i/_0500_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0803_  (.A(net679),
    .B(\i_ibex/lsu_addr_last [24]),
    .X(\i_ibex/id_stage_i/_0502_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0804_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net352),
    .C1(\i_ibex/id_stage_i/_0502_ ),
    .B1(\i_ibex/id_stage_i/_0368_ ),
    .A1(\i_ibex/pc_id [24]),
    .Y(\i_ibex/id_stage_i/_0503_ ),
    .A2(\i_ibex/id_stage_i/_0366_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0805_  (.B1(\i_ibex/id_stage_i/_0503_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [24]),
    .VSS(VSS),
    .A1(net1304),
    .A2(\i_ibex/id_stage_i/_0501_ ));
 sg13g2_and3_2 \i_ibex/id_stage_i/_0806_  (.X(\i_ibex/id_stage_i/_0504_ ),
    .A(net1380),
    .B(net1261),
    .C(\i_ibex/rf_rdata_a [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0807_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1297),
    .A2(\i_ibex/lsu_addr_last [23]),
    .Y(\i_ibex/id_stage_i/_0505_ ),
    .B1(\i_ibex/id_stage_i/_0504_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0808_  (.A(net679),
    .B(\i_ibex/lsu_addr_last [23]),
    .X(\i_ibex/id_stage_i/_0506_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0809_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net353),
    .C1(\i_ibex/id_stage_i/_0506_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [23]),
    .Y(\i_ibex/id_stage_i/_0507_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0810_  (.B1(\i_ibex/id_stage_i/_0507_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [23]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0505_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0811_  (.X(\i_ibex/id_stage_i/_0508_ ),
    .A(net1378),
    .B(net1259),
    .C(\i_ibex/rf_rdata_a [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0812_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1299),
    .A2(\i_ibex/lsu_addr_last [22]),
    .Y(\i_ibex/id_stage_i/_0509_ ),
    .B1(\i_ibex/id_stage_i/_0508_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0813_  (.A(net679),
    .B(\i_ibex/lsu_addr_last [22]),
    .X(\i_ibex/id_stage_i/_0510_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0814_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net354),
    .C1(\i_ibex/id_stage_i/_0510_ ),
    .B1(net1196),
    .A1(\i_ibex/pc_id [22]),
    .Y(\i_ibex/id_stage_i/_0511_ ),
    .A2(net1257));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_0815_  (.B1(\i_ibex/id_stage_i/_0511_ ),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_a_ex [22]),
    .VSS(VSS),
    .A1(net1302),
    .A2(\i_ibex/id_stage_i/_0509_ ));
 sg13g2_buf_2 fanout668 (.A(net672),
    .X(net668),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout667 (.A(net672),
    .X(net667),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0818_  (.Y(\i_ibex/id_stage_i/_0514_ ),
    .B(\i_ibex/rf_rdata_b [31]),
    .A_N(net1366),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout666 (.A(\i_ibex/if_stage_i/fetch_rdata [14]),
    .X(net666),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout665 (.A(\i_ibex/if_stage_i/fetch_rdata [14]),
    .X(net665),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0821_  (.A0(net722),
    .A1(net722),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0517_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_0822_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0518_ ),
    .A(net1329),
    .VSS(VSS));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_0824_  (.X(\i_ibex/id_stage_i/_0520_ ),
    .A(net1381),
    .B(\i_ibex/id_stage_i/_0518_ ),
    .C(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout663 (.A(net666),
    .X(net663),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/_0826_  (.A(net679),
    .B(net1328),
    .C(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .Y(\i_ibex/id_stage_i/_0522_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_0827_  (.A(net677),
    .B(\i_ibex/id_stage_i/_0522_ ),
    .X(\i_ibex/id_stage_i/_0523_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(net666),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout661 (.A(net665),
    .X(net661),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout660 (.A(net665),
    .X(net660),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0831_  (.Y(\i_ibex/id_stage_i/_0527_ ),
    .B(net722),
    .A_N(net1327),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout659 (.A(net665),
    .X(net659),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0833_  (.Y(\i_ibex/id_stage_i/_0529_ ),
    .A(net1327),
    .B(net722),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/id_stage_i/_0834_  (.A(net688),
    .B(net678),
    .C(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .X(\i_ibex/id_stage_i/_0530_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout658 (.A(net665),
    .X(net658),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0836_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0527_ ),
    .A2(\i_ibex/id_stage_i/_0529_ ),
    .Y(\i_ibex/id_stage_i/_0532_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0837_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net722),
    .C1(\i_ibex/id_stage_i/_0532_ ),
    .B1(net1188),
    .A1(\i_ibex/id_stage_i/_0517_ ),
    .Y(\i_ibex/id_stage_i/_0533_ ),
    .A2(net1249));
 sg13g2_buf_2 fanout657 (.A(\i_ibex/if_stage_i/fetch_rdata [13]),
    .X(net657),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout656 (.A(net657),
    .X(net656),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout655 (.A(net657),
    .X(net655),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0841_  (.Y(\i_ibex/id_stage_i/_0537_ ),
    .A(net1331),
    .B(net677),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net657),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0843_  (.B(net1368),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0539_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0533_ ));
 sg13g2_buf_2 fanout653 (.A(net657),
    .X(net653),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0845_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [31]),
    .A2(\i_ibex/id_stage_i/_0539_ ),
    .A1(\i_ibex/id_stage_i/_0514_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0846_  (.Y(\i_ibex/id_stage_i/_0541_ ),
    .B(\i_ibex/rf_rdata_b [30]),
    .A_N(net1369),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0847_  (.A0(net722),
    .A1(net734),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0542_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout652 (.A(net657),
    .X(net652),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0849_  (.Y(\i_ibex/id_stage_i/_0544_ ),
    .B(net722),
    .A_N(net1328),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0850_  (.Y(\i_ibex/id_stage_i/_0545_ ),
    .A(net1328),
    .B(net722),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0851_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0544_ ),
    .A2(\i_ibex/id_stage_i/_0545_ ),
    .Y(\i_ibex/id_stage_i/_0546_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0852_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0546_ ),
    .B1(\i_ibex/id_stage_i/_0542_ ),
    .A1(net723),
    .Y(\i_ibex/id_stage_i/_0547_ ),
    .A2(net1188));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0853_  (.B(net1369),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0548_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0547_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0854_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [30]),
    .A2(\i_ibex/id_stage_i/_0548_ ),
    .A1(\i_ibex/id_stage_i/_0541_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0855_  (.Y(\i_ibex/id_stage_i/_0549_ ),
    .B(\i_ibex/rf_rdata_b [21]),
    .A_N(net1370),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0856_  (.A0(net723),
    .A1(net757),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0550_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0857_  (.Y(\i_ibex/id_stage_i/_0551_ ),
    .B(net723),
    .A_N(net1328),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0858_  (.Y(\i_ibex/id_stage_i/_0552_ ),
    .A(net1328),
    .B(net723),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0859_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0551_ ),
    .A2(\i_ibex/id_stage_i/_0552_ ),
    .Y(\i_ibex/id_stage_i/_0553_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0860_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0553_ ),
    .B1(\i_ibex/id_stage_i/_0550_ ),
    .A1(net723),
    .Y(\i_ibex/id_stage_i/_0554_ ),
    .A2(net1188));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0861_  (.B(net1369),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0555_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0554_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0862_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [21]),
    .A2(\i_ibex/id_stage_i/_0555_ ),
    .A1(\i_ibex/id_stage_i/_0549_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0863_  (.Y(\i_ibex/id_stage_i/_0556_ ),
    .B(\i_ibex/rf_rdata_b [20]),
    .A_N(net1369),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0864_  (.A0(net723),
    .A1(net761),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0557_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0865_  (.Y(\i_ibex/id_stage_i/_0558_ ),
    .B(net723),
    .A_N(net1333),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0866_  (.Y(\i_ibex/id_stage_i/_0069_ ),
    .A(net1333),
    .B(net723),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0867_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0558_ ),
    .A2(\i_ibex/id_stage_i/_0069_ ),
    .Y(\i_ibex/id_stage_i/_0070_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0868_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0070_ ),
    .B1(\i_ibex/id_stage_i/_0557_ ),
    .A1(net724),
    .Y(\i_ibex/id_stage_i/_0071_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0869_  (.B(net1369),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0072_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0071_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0870_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [20]),
    .A2(\i_ibex/id_stage_i/_0072_ ),
    .A1(\i_ibex/id_stage_i/_0556_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0871_  (.Y(\i_ibex/id_stage_i/_0073_ ),
    .B(\i_ibex/rf_rdata_b [19]),
    .A_N(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0872_  (.A0(net724),
    .A1(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0873_  (.Y(\i_ibex/id_stage_i/_0075_ ),
    .B(net724),
    .A_N(net1333),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0874_  (.Y(\i_ibex/id_stage_i/_0076_ ),
    .A(net1333),
    .B(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0875_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0075_ ),
    .A2(\i_ibex/id_stage_i/_0076_ ),
    .Y(\i_ibex/id_stage_i/_0077_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0876_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0077_ ),
    .B1(\i_ibex/id_stage_i/_0074_ ),
    .A1(net724),
    .Y(\i_ibex/id_stage_i/_0078_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0877_  (.B(net1375),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0078_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0878_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net683),
    .Y(\i_ibex/alu_operand_b_ex [19]),
    .A2(\i_ibex/id_stage_i/_0079_ ),
    .A1(\i_ibex/id_stage_i/_0073_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0879_  (.Y(\i_ibex/id_stage_i/_0080_ ),
    .B(\i_ibex/rf_rdata_b [18]),
    .A_N(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0880_  (.A0(net724),
    .A1(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout651 (.A(net657),
    .X(net651),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0882_  (.Y(\i_ibex/id_stage_i/_0083_ ),
    .B(net724),
    .A_N(net1332),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0883_  (.Y(\i_ibex/id_stage_i/_0084_ ),
    .A(net1332),
    .B(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0884_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0083_ ),
    .A2(\i_ibex/id_stage_i/_0084_ ),
    .Y(\i_ibex/id_stage_i/_0085_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0885_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0085_ ),
    .B1(\i_ibex/id_stage_i/_0081_ ),
    .A1(net724),
    .Y(\i_ibex/id_stage_i/_0086_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0886_  (.B(net1375),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0087_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0086_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0887_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net683),
    .Y(\i_ibex/alu_operand_b_ex [18]),
    .A2(\i_ibex/id_stage_i/_0087_ ),
    .A1(\i_ibex/id_stage_i/_0080_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0888_  (.Y(\i_ibex/id_stage_i/_0088_ ),
    .B(\i_ibex/rf_rdata_b [17]),
    .A_N(net1374),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0889_  (.A0(net724),
    .A1(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0089_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0890_  (.Y(\i_ibex/id_stage_i/_0090_ ),
    .B(net725),
    .A_N(net1333),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0891_  (.Y(\i_ibex/id_stage_i/_0091_ ),
    .A(net1337),
    .B(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0892_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0090_ ),
    .A2(\i_ibex/id_stage_i/_0091_ ),
    .Y(\i_ibex/id_stage_i/_0092_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0893_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0092_ ),
    .B1(\i_ibex/id_stage_i/_0089_ ),
    .A1(net725),
    .Y(\i_ibex/id_stage_i/_0093_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0894_  (.B(net1375),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0094_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0093_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0895_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net683),
    .Y(\i_ibex/alu_operand_b_ex [17]),
    .A2(\i_ibex/id_stage_i/_0094_ ),
    .A1(\i_ibex/id_stage_i/_0088_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0896_  (.Y(\i_ibex/id_stage_i/_0095_ ),
    .B(\i_ibex/rf_rdata_b [16]),
    .A_N(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout650 (.A(net657),
    .X(net650),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0898_  (.A0(net725),
    .A1(net766),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0899_  (.Y(\i_ibex/id_stage_i/_0098_ ),
    .A(net1334),
    .B(net766),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0900_  (.Y(\i_ibex/id_stage_i/_0099_ ),
    .B(net725),
    .A_N(net1334),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0901_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0098_ ),
    .A2(\i_ibex/id_stage_i/_0099_ ),
    .Y(\i_ibex/id_stage_i/_0100_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0902_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0100_ ),
    .B1(\i_ibex/id_stage_i/_0097_ ),
    .A1(net725),
    .Y(\i_ibex/id_stage_i/_0101_ ),
    .A2(net1191));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0903_  (.B(net1374),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0102_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0101_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0904_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net683),
    .Y(\i_ibex/alu_operand_b_ex [16]),
    .A2(\i_ibex/id_stage_i/_0102_ ),
    .A1(\i_ibex/id_stage_i/_0095_ ));
 sg13g2_buf_2 fanout649 (.A(\i_ibex/if_stage_i/fetch_rdata [12]),
    .X(net649),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0906_  (.Y(\i_ibex/id_stage_i/_0104_ ),
    .B(\i_ibex/rf_rdata_b [15]),
    .A_N(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0907_  (.A0(net725),
    .A1(net768),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0908_  (.Y(\i_ibex/id_stage_i/_0106_ ),
    .A(net1335),
    .B(net768),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0909_  (.Y(\i_ibex/id_stage_i/_0107_ ),
    .B(net725),
    .A_N(net1335),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0910_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0106_ ),
    .A2(\i_ibex/id_stage_i/_0107_ ),
    .Y(\i_ibex/id_stage_i/_0108_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0911_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0108_ ),
    .B1(\i_ibex/id_stage_i/_0105_ ),
    .A1(net725),
    .Y(\i_ibex/id_stage_i/_0109_ ),
    .A2(net1191));
 sg13g2_buf_2 fanout648 (.A(\i_ibex/if_stage_i/fetch_rdata [12]),
    .X(net648),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0913_  (.B(net1375),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0111_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0109_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0914_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net683),
    .Y(\i_ibex/alu_operand_b_ex [15]),
    .A2(\i_ibex/id_stage_i/_0111_ ),
    .A1(\i_ibex/id_stage_i/_0104_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0915_  (.Y(\i_ibex/id_stage_i/_0112_ ),
    .B(\i_ibex/rf_rdata_b [14]),
    .A_N(net1372),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0916_  (.A0(net726),
    .A1(net770),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0917_  (.Y(\i_ibex/id_stage_i/_0114_ ),
    .A(net1334),
    .B(net770),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0918_  (.Y(\i_ibex/id_stage_i/_0115_ ),
    .B(net726),
    .A_N(net1335),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0919_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0114_ ),
    .A2(\i_ibex/id_stage_i/_0115_ ),
    .Y(\i_ibex/id_stage_i/_0116_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0920_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0116_ ),
    .B1(\i_ibex/id_stage_i/_0113_ ),
    .A1(net726),
    .Y(\i_ibex/id_stage_i/_0117_ ),
    .A2(net1191));
 sg13g2_buf_2 fanout647 (.A(\i_ibex/if_stage_i/fetch_rdata [12]),
    .X(net647),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0922_  (.B(net1372),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0119_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0117_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0923_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net683),
    .Y(\i_ibex/alu_operand_b_ex [14]),
    .A2(\i_ibex/id_stage_i/_0119_ ),
    .A1(\i_ibex/id_stage_i/_0112_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0924_  (.Y(\i_ibex/id_stage_i/_0120_ ),
    .B(\i_ibex/rf_rdata_b [13]),
    .A_N(net1374),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout646 (.A(\i_ibex/if_stage_i/fetch_rdata [12]),
    .X(net646),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0926_  (.A0(net726),
    .A1(net774),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0927_  (.Y(\i_ibex/id_stage_i/_0123_ ),
    .A(net1334),
    .B(net774),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0928_  (.Y(\i_ibex/id_stage_i/_0124_ ),
    .B(net726),
    .A_N(net1335),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout645 (.A(\i_ibex/if_stage_i/fetch_rdata [11]),
    .X(net645),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0930_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0123_ ),
    .A2(\i_ibex/id_stage_i/_0124_ ),
    .Y(\i_ibex/id_stage_i/_0126_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0931_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0126_ ),
    .B1(\i_ibex/id_stage_i/_0122_ ),
    .A1(net726),
    .Y(\i_ibex/id_stage_i/_0127_ ),
    .A2(net1191));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0932_  (.B(net1374),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0127_ ));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(\i_ibex/if_stage_i/fetch_rdata [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0934_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [13]),
    .A2(\i_ibex/id_stage_i/_0128_ ),
    .A1(\i_ibex/id_stage_i/_0120_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0935_  (.Y(\i_ibex/id_stage_i/_0130_ ),
    .B(\i_ibex/rf_rdata_b [12]),
    .A_N(net1372),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0936_  (.A0(net726),
    .A1(net778),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout643 (.A(\i_ibex/if_stage_i/fetch_rdata [8]),
    .X(net643),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0938_  (.Y(\i_ibex/id_stage_i/_0133_ ),
    .A(net1336),
    .B(net778),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0939_  (.Y(\i_ibex/id_stage_i/_0134_ ),
    .B(net726),
    .A_N(net1336),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0940_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0133_ ),
    .A2(\i_ibex/id_stage_i/_0134_ ),
    .Y(\i_ibex/id_stage_i/_0135_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0941_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0135_ ),
    .B1(\i_ibex/id_stage_i/_0131_ ),
    .A1(net727),
    .Y(\i_ibex/id_stage_i/_0136_ ),
    .A2(net1191));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0942_  (.B(net1372),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0137_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0136_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0943_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [12]),
    .A2(\i_ibex/id_stage_i/_0137_ ),
    .A1(\i_ibex/id_stage_i/_0130_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0944_  (.Y(\i_ibex/id_stage_i/_0138_ ),
    .B(\i_ibex/rf_rdata_b [29]),
    .A_N(net1373),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0945_  (.A0(net727),
    .A1(net741),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0139_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(\i_ibex/if_stage_i/fetch_rdata [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0947_  (.Y(\i_ibex/id_stage_i/_0141_ ),
    .A(net1336),
    .B(net727),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0948_  (.Y(\i_ibex/id_stage_i/_0142_ ),
    .B(net727),
    .A_N(net1336),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0949_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0141_ ),
    .A2(\i_ibex/id_stage_i/_0142_ ),
    .Y(\i_ibex/id_stage_i/_0143_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0950_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0143_ ),
    .B1(\i_ibex/id_stage_i/_0139_ ),
    .A1(net727),
    .Y(\i_ibex/id_stage_i/_0144_ ),
    .A2(net1191));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0951_  (.B(net1372),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0145_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0144_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0952_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [29]),
    .A2(\i_ibex/id_stage_i/_0145_ ),
    .A1(\i_ibex/id_stage_i/_0138_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0953_  (.Y(\i_ibex/id_stage_i/_0146_ ),
    .B(\i_ibex/rf_rdata_b [11]),
    .A_N(net1366),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0954_  (.A0(net727),
    .A1(net355),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0955_  (.Y(\i_ibex/id_stage_i/_0148_ ),
    .A(net1328),
    .B(net761),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0956_  (.Y(\i_ibex/id_stage_i/_0149_ ),
    .B(net727),
    .A_N(net1327),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0957_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0148_ ),
    .A2(\i_ibex/id_stage_i/_0149_ ),
    .Y(\i_ibex/id_stage_i/_0150_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0958_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1250),
    .C1(\i_ibex/id_stage_i/_0150_ ),
    .B1(\i_ibex/id_stage_i/_0147_ ),
    .A1(\i_ibex/id_stage_i/imm_s_type [0]),
    .Y(\i_ibex/id_stage_i/_0151_ ),
    .A2(net1189));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0959_  (.B(net1367),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0152_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0151_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0960_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [11]),
    .A2(\i_ibex/id_stage_i/_0152_ ),
    .A1(\i_ibex/id_stage_i/_0146_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0961_  (.Y(\i_ibex/id_stage_i/_0153_ ),
    .B(\i_ibex/rf_rdata_b [10]),
    .A_N(net1366),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0962_  (.A0(net734),
    .A1(net356),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0963_  (.Y(\i_ibex/id_stage_i/_0155_ ),
    .A(net1327),
    .B(net734),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0964_  (.Y(\i_ibex/id_stage_i/_0156_ ),
    .B(net734),
    .A_N(net1327),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0965_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0155_ ),
    .A2(\i_ibex/id_stage_i/_0156_ ),
    .Y(\i_ibex/id_stage_i/_0157_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0966_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0157_ ),
    .B1(\i_ibex/id_stage_i/_0154_ ),
    .A1(net734),
    .Y(\i_ibex/id_stage_i/_0158_ ),
    .A2(net1188));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0967_  (.B(net1367),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0158_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0968_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [10]),
    .A2(\i_ibex/id_stage_i/_0159_ ),
    .A1(\i_ibex/id_stage_i/_0153_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0969_  (.Y(\i_ibex/id_stage_i/_0160_ ),
    .B(\i_ibex/rf_rdata_b [9]),
    .A_N(net1370),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0970_  (.A0(net741),
    .A1(net357),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0971_  (.Y(\i_ibex/id_stage_i/_0162_ ),
    .A(net1333),
    .B(net741),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(\i_ibex/if_stage_i/fetch_rdata [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0973_  (.Y(\i_ibex/id_stage_i/_0164_ ),
    .B(net741),
    .A_N(net1333),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0974_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0162_ ),
    .A2(\i_ibex/id_stage_i/_0164_ ),
    .Y(\i_ibex/id_stage_i/_0165_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0975_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0165_ ),
    .B1(\i_ibex/id_stage_i/_0161_ ),
    .A1(net742),
    .Y(\i_ibex/id_stage_i/_0166_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0976_  (.B(net1372),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0167_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0166_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0977_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [9]),
    .A2(\i_ibex/id_stage_i/_0167_ ),
    .A1(\i_ibex/id_stage_i/_0160_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0978_  (.Y(\i_ibex/id_stage_i/_0168_ ),
    .B(\i_ibex/rf_rdata_b [8]),
    .A_N(net1370),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0979_  (.A0(net743),
    .A1(net358),
    .S(net674),
    .X(\i_ibex/id_stage_i/_0169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0980_  (.Y(\i_ibex/id_stage_i/_0170_ ),
    .A(net1329),
    .B(net743),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0981_  (.Y(\i_ibex/id_stage_i/_0171_ ),
    .B(net743),
    .A_N(net1331),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0982_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0170_ ),
    .A2(\i_ibex/id_stage_i/_0171_ ),
    .Y(\i_ibex/id_stage_i/_0172_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0983_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0172_ ),
    .B1(\i_ibex/id_stage_i/_0169_ ),
    .A1(net744),
    .Y(\i_ibex/id_stage_i/_0173_ ),
    .A2(net1188));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0984_  (.B(net1369),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0174_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0173_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0985_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [8]),
    .A2(\i_ibex/id_stage_i/_0174_ ),
    .A1(\i_ibex/id_stage_i/_0168_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0986_  (.Y(\i_ibex/id_stage_i/_0175_ ),
    .B(\i_ibex/rf_rdata_b [7]),
    .A_N(net1367),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout640 (.A(\i_ibex/if_stage_i/fetch_rdata [0]),
    .X(net640),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0988_  (.A0(net745),
    .A1(net359),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0177_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0989_  (.Y(\i_ibex/id_stage_i/_0178_ ),
    .A(net1330),
    .B(net745),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0990_  (.Y(\i_ibex/id_stage_i/_0179_ ),
    .B(net745),
    .A_N(net1330),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_0991_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0178_ ),
    .A2(\i_ibex/id_stage_i/_0179_ ),
    .Y(\i_ibex/id_stage_i/_0180_ ),
    .B1(net1245));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_0992_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1250),
    .C1(\i_ibex/id_stage_i/_0180_ ),
    .B1(\i_ibex/id_stage_i/_0177_ ),
    .A1(net746),
    .Y(\i_ibex/id_stage_i/_0181_ ),
    .A2(net1189));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_0993_  (.B(net1367),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0182_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0181_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_0994_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [7]),
    .A2(\i_ibex/id_stage_i/_0182_ ),
    .A1(\i_ibex/id_stage_i/_0175_ ));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0996_  (.Y(\i_ibex/id_stage_i/_0184_ ),
    .B(\i_ibex/rf_rdata_b [6]),
    .A_N(net1366),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_0997_  (.A0(net747),
    .A1(net360),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_0998_  (.Y(\i_ibex/id_stage_i/_0186_ ),
    .A(net1330),
    .B(net747),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_0999_  (.Y(\i_ibex/id_stage_i/_0187_ ),
    .B(net747),
    .A_N(net1330),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1000_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0186_ ),
    .A2(\i_ibex/id_stage_i/_0187_ ),
    .Y(\i_ibex/id_stage_i/_0188_ ),
    .B1(net1245));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1001_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1250),
    .C1(\i_ibex/id_stage_i/_0188_ ),
    .B1(\i_ibex/id_stage_i/_0185_ ),
    .A1(net747),
    .Y(\i_ibex/id_stage_i/_0189_ ),
    .A2(net1188));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(net640),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1003_  (.B(net1366),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0191_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0189_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1004_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [6]),
    .A2(\i_ibex/id_stage_i/_0191_ ),
    .A1(\i_ibex/id_stage_i/_0184_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1005_  (.Y(\i_ibex/id_stage_i/_0192_ ),
    .B(\i_ibex/rf_rdata_b [5]),
    .A_N(net1368),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1006_  (.A0(net750),
    .A1(net361),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1007_  (.Y(\i_ibex/id_stage_i/_0194_ ),
    .A(net1329),
    .B(net750),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1008_  (.Y(\i_ibex/id_stage_i/_0195_ ),
    .B(net750),
    .A_N(net1331),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1009_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0194_ ),
    .A2(\i_ibex/id_stage_i/_0195_ ),
    .Y(\i_ibex/id_stage_i/_0196_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1010_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1250),
    .C1(\i_ibex/id_stage_i/_0196_ ),
    .B1(\i_ibex/id_stage_i/_0193_ ),
    .A1(net752),
    .Y(\i_ibex/id_stage_i/_0197_ ),
    .A2(net1188));
 sg13g2_buf_2 fanout637 (.A(net640),
    .X(net637),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1012_  (.B(net1369),
    .C(\i_ibex/id_stage_i/_0537_ ),
    .Y(\i_ibex/id_stage_i/_0199_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0197_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1013_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net684),
    .Y(\i_ibex/alu_operand_b_ex [5]),
    .A2(\i_ibex/id_stage_i/_0199_ ),
    .A1(\i_ibex/id_stage_i/_0192_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1014_  (.Y(\i_ibex/id_stage_i/_0200_ ),
    .B(\i_ibex/rf_rdata_b [4]),
    .A_N(net1367),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout636 (.A(net640),
    .X(net636),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1016_  (.A0(\i_ibex/id_stage_i/imm_s_type [4]),
    .A1(net362),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1017_  (.Y(\i_ibex/id_stage_i/_0203_ ),
    .A(net1330),
    .B(net753),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1018_  (.Y(\i_ibex/id_stage_i/_0204_ ),
    .B(net753),
    .A_N(net1330),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout635 (.A(\i_ibex/load_store_unit_i/_0236_ ),
    .X(net635),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1020_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0203_ ),
    .A2(\i_ibex/id_stage_i/_0204_ ),
    .Y(\i_ibex/id_stage_i/_0206_ ),
    .B1(net1245));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1021_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1250),
    .C1(\i_ibex/id_stage_i/_0206_ ),
    .B1(\i_ibex/id_stage_i/_0202_ ),
    .A1(\i_ibex/id_stage_i/imm_s_type [4]),
    .Y(\i_ibex/id_stage_i/_0207_ ),
    .A2(net1189));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1022_  (.B(net1371),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0208_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0207_ ));
 sg13g2_buf_2 fanout634 (.A(\i_ibex/cs_registers_i/_0150_ ),
    .X(net634),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1024_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [4]),
    .A2(\i_ibex/id_stage_i/_0208_ ),
    .A1(\i_ibex/id_stage_i/_0200_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1025_  (.Y(\i_ibex/id_stage_i/_0210_ ),
    .B(\i_ibex/rf_rdata_b [3]),
    .A_N(net1366),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1026_  (.A0(\i_ibex/id_stage_i/imm_s_type [3]),
    .A1(net363),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1027_  (.Y(\i_ibex/id_stage_i/_0212_ ),
    .A(net1330),
    .B(net754),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1028_  (.Y(\i_ibex/id_stage_i/_0213_ ),
    .B(net754),
    .A_N(net1330),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1029_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0212_ ),
    .A2(\i_ibex/id_stage_i/_0213_ ),
    .Y(\i_ibex/id_stage_i/_0214_ ),
    .B1(net1245));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1030_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1250),
    .C1(\i_ibex/id_stage_i/_0214_ ),
    .B1(\i_ibex/id_stage_i/_0211_ ),
    .A1(\i_ibex/id_stage_i/imm_s_type [3]),
    .Y(\i_ibex/id_stage_i/_0215_ ),
    .A2(net1189));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1031_  (.B(net1366),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0216_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0215_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1032_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [3]),
    .A2(\i_ibex/id_stage_i/_0216_ ),
    .A1(\i_ibex/id_stage_i/_0210_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/_1033_  (.A(net1366),
    .B(\i_ibex/rf_rdata_b [2]),
    .Y(\i_ibex/id_stage_i/_0217_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1034_  (.Y(\i_ibex/id_stage_i/_0218_ ),
    .A(\i_ibex/id_stage_i/imm_b_mux_sel_dec [1]),
    .B(net364),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1035_  (.Y(\i_ibex/id_stage_i/_0219_ ),
    .B(\i_ibex/id_stage_i/imm_s_type [2]),
    .A_N(net677),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1036_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0218_ ),
    .A2(\i_ibex/id_stage_i/_0219_ ),
    .Y(\i_ibex/id_stage_i/_0220_ ),
    .B1(net1329));
 sg13g2_nor3_1 \i_ibex/id_stage_i/_1037_  (.A(\i_ibex/id_stage_i/_0518_ ),
    .B(\i_ibex/id_stage_i/imm_b_mux_sel_dec [1]),
    .C(net783),
    .Y(\i_ibex/id_stage_i/_0221_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1038_  (.B1(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0222_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/_0220_ ),
    .A2(\i_ibex/id_stage_i/_0221_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/_1039_  (.A(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .B_N(net755),
    .Y(\i_ibex/id_stage_i/_0223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1040_  (.B1(net1329),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0224_ ),
    .VSS(VSS),
    .A1(net677),
    .A2(\i_ibex/id_stage_i/_0223_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/_1041_  (.A(net678),
    .B_N(net755),
    .Y(\i_ibex/id_stage_i/_0225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/_1042_  (.Y(\i_ibex/id_stage_i/_0226_ ),
    .B1(\i_ibex/id_stage_i/_0225_ ),
    .B2(\i_ibex/id_stage_i/_0518_ ),
    .A2(\i_ibex/id_stage_i/imm_s_type [2]),
    .A1(net678),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/_1043_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/_0227_ ),
    .B(\i_ibex/id_stage_i/_0226_ ),
    .A(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]));
 sg13g2_and4_1 \i_ibex/id_stage_i/_1044_  (.A(net1371),
    .B(\i_ibex/id_stage_i/_0222_ ),
    .C(\i_ibex/id_stage_i/_0224_ ),
    .D(\i_ibex/id_stage_i/_0227_ ),
    .X(\i_ibex/id_stage_i/_0228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1045_  (.B1(net1381),
    .VDD(VDD),
    .Y(\i_ibex/alu_operand_b_ex [2]),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/_0217_ ),
    .A2(\i_ibex/id_stage_i/_0228_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1046_  (.Y(\i_ibex/id_stage_i/_0229_ ),
    .B(\i_ibex/rf_rdata_b [28]),
    .A_N(net1369),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1047_  (.A0(net727),
    .A1(net743),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0230_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1048_  (.Y(\i_ibex/id_stage_i/_0231_ ),
    .A(net1329),
    .B(net728),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1049_  (.Y(\i_ibex/id_stage_i/_0232_ ),
    .B(net728),
    .A_N(net1329),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1050_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0231_ ),
    .A2(\i_ibex/id_stage_i/_0232_ ),
    .Y(\i_ibex/id_stage_i/_0233_ ),
    .B1(net1245));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1051_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0233_ ),
    .B1(\i_ibex/id_stage_i/_0230_ ),
    .A1(net728),
    .Y(\i_ibex/id_stage_i/_0234_ ),
    .A2(net1189));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1052_  (.B(net1370),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0235_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0234_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1053_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [28]),
    .A2(\i_ibex/id_stage_i/_0235_ ),
    .A1(\i_ibex/id_stage_i/_0229_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1054_  (.Y(\i_ibex/id_stage_i/_0236_ ),
    .B(\i_ibex/rf_rdata_b [1]),
    .A_N(net1368),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1055_  (.A0(net757),
    .A1(\i_ibex/id_stage_i/imm_s_type [1]),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1056_  (.Y(\i_ibex/id_stage_i/_0238_ ),
    .A(\i_ibex/id_stage_i/_0522_ ),
    .B(\i_ibex/id_stage_i/_0237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1057_  (.A0(net757),
    .A1(net783),
    .S(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .X(\i_ibex/id_stage_i/_0239_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1058_  (.A0(\i_ibex/id_stage_i/imm_s_type [1]),
    .A1(net365),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0240_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/_1059_  (.A(net1327),
    .B_N(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .Y(\i_ibex/id_stage_i/_0241_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/_1060_  (.Y(\i_ibex/id_stage_i/_0242_ ),
    .B1(\i_ibex/id_stage_i/_0240_ ),
    .B2(\i_ibex/id_stage_i/_0241_ ),
    .A2(\i_ibex/id_stage_i/_0239_ ),
    .A1(net1327),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1061_  (.Y(\i_ibex/id_stage_i/_0243_ ),
    .A(\i_ibex/id_stage_i/_0238_ ),
    .B(\i_ibex/id_stage_i/_0242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/_1062_  (.B(net1240),
    .C(\i_ibex/id_stage_i/_0243_ ),
    .A(net1367),
    .Y(\i_ibex/id_stage_i/_0244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1063_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [1]),
    .A2(\i_ibex/id_stage_i/_0244_ ),
    .A1(\i_ibex/id_stage_i/_0236_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1064_  (.Y(\i_ibex/id_stage_i/_0245_ ),
    .B(\i_ibex/rf_rdata_b [0]),
    .A_N(net1367),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1065_  (.A0(\i_ibex/id_stage_i/imm_s_type [0]),
    .A1(net366),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0246_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1066_  (.Y(\i_ibex/id_stage_i/_0247_ ),
    .A(net1327),
    .B(net367),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1067_  (.Y(\i_ibex/id_stage_i/_0248_ ),
    .B(net761),
    .A_N(net1328),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1068_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0247_ ),
    .A2(\i_ibex/id_stage_i/_0248_ ),
    .Y(\i_ibex/id_stage_i/_0249_ ),
    .B1(net1244));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1069_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0249_ ),
    .B1(\i_ibex/id_stage_i/_0246_ ),
    .A1(net368),
    .Y(\i_ibex/id_stage_i/_0250_ ),
    .A2(net1188));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1070_  (.B(net1367),
    .C(net1240),
    .Y(\i_ibex/id_stage_i/_0251_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0250_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1071_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0245_ ),
    .A2(\i_ibex/id_stage_i/_0251_ ),
    .Y(\i_ibex/alu_operand_b_ex [0]),
    .B1(net686));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1072_  (.Y(\i_ibex/id_stage_i/_0252_ ),
    .B(\i_ibex/rf_rdata_b [27]),
    .A_N(net1370),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1073_  (.A0(net728),
    .A1(net745),
    .S(net676),
    .X(\i_ibex/id_stage_i/_0253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1074_  (.Y(\i_ibex/id_stage_i/_0254_ ),
    .A(net1329),
    .B(net728),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1075_  (.Y(\i_ibex/id_stage_i/_0255_ ),
    .B(net728),
    .A_N(net1331),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1076_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0254_ ),
    .A2(\i_ibex/id_stage_i/_0255_ ),
    .Y(\i_ibex/id_stage_i/_0256_ ),
    .B1(net1245));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1077_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1249),
    .C1(\i_ibex/id_stage_i/_0256_ ),
    .B1(\i_ibex/id_stage_i/_0253_ ),
    .A1(net728),
    .Y(\i_ibex/id_stage_i/_0257_ ),
    .A2(net1189));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1078_  (.B(net1370),
    .C(net1241),
    .Y(\i_ibex/id_stage_i/_0258_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0257_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1079_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [27]),
    .A2(\i_ibex/id_stage_i/_0258_ ),
    .A1(\i_ibex/id_stage_i/_0252_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1080_  (.Y(\i_ibex/id_stage_i/_0259_ ),
    .B(\i_ibex/rf_rdata_b [26]),
    .A_N(net1373),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1081_  (.A0(net728),
    .A1(net747),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1082_  (.Y(\i_ibex/id_stage_i/_0261_ ),
    .A(net1334),
    .B(net729),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1083_  (.Y(\i_ibex/id_stage_i/_0262_ ),
    .B(net729),
    .A_N(net1334),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1084_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0261_ ),
    .A2(\i_ibex/id_stage_i/_0262_ ),
    .Y(\i_ibex/id_stage_i/_0263_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1085_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0263_ ),
    .B1(\i_ibex/id_stage_i/_0260_ ),
    .A1(net729),
    .Y(\i_ibex/id_stage_i/_0264_ ),
    .A2(net1191));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1086_  (.B(net1373),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0265_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0264_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1087_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [26]),
    .A2(\i_ibex/id_stage_i/_0265_ ),
    .A1(\i_ibex/id_stage_i/_0259_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1088_  (.Y(\i_ibex/id_stage_i/_0266_ ),
    .B(\i_ibex/rf_rdata_b [25]),
    .A_N(net1372),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1089_  (.A0(net729),
    .A1(net750),
    .S(net675),
    .X(\i_ibex/id_stage_i/_0267_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1090_  (.Y(\i_ibex/id_stage_i/_0268_ ),
    .A(net1334),
    .B(net729),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1091_  (.Y(\i_ibex/id_stage_i/_0269_ ),
    .B(net729),
    .A_N(net1334),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1092_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0268_ ),
    .A2(\i_ibex/id_stage_i/_0269_ ),
    .Y(\i_ibex/id_stage_i/_0270_ ),
    .B1(net1247));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1093_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1252),
    .C1(\i_ibex/id_stage_i/_0270_ ),
    .B1(\i_ibex/id_stage_i/_0267_ ),
    .A1(net729),
    .Y(\i_ibex/id_stage_i/_0271_ ),
    .A2(net1191));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1094_  (.B(net1372),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0272_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0271_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1095_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net686),
    .Y(\i_ibex/alu_operand_b_ex [25]),
    .A2(\i_ibex/id_stage_i/_0272_ ),
    .A1(\i_ibex/id_stage_i/_0266_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1096_  (.Y(\i_ibex/id_stage_i/_0273_ ),
    .B(\i_ibex/rf_rdata_b [24]),
    .A_N(net1374),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1097_  (.A0(net729),
    .A1(net753),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1098_  (.Y(\i_ibex/id_stage_i/_0275_ ),
    .A(net1332),
    .B(net730),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1099_  (.Y(\i_ibex/id_stage_i/_0276_ ),
    .B(net730),
    .A_N(net1332),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1100_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0275_ ),
    .A2(\i_ibex/id_stage_i/_0276_ ),
    .Y(\i_ibex/id_stage_i/_0277_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1101_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0277_ ),
    .B1(\i_ibex/id_stage_i/_0274_ ),
    .A1(net730),
    .Y(\i_ibex/id_stage_i/_0278_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1102_  (.B(net1374),
    .C(net1243),
    .Y(\i_ibex/id_stage_i/_0279_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0278_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1103_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [24]),
    .A2(\i_ibex/id_stage_i/_0279_ ),
    .A1(\i_ibex/id_stage_i/_0273_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1104_  (.Y(\i_ibex/id_stage_i/_0280_ ),
    .B(\i_ibex/rf_rdata_b [23]),
    .A_N(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1105_  (.A0(net730),
    .A1(net754),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0281_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1106_  (.Y(\i_ibex/id_stage_i/_0282_ ),
    .A(net1332),
    .B(net730),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1107_  (.Y(\i_ibex/id_stage_i/_0283_ ),
    .B(net730),
    .A_N(net1332),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1108_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0282_ ),
    .A2(\i_ibex/id_stage_i/_0283_ ),
    .Y(\i_ibex/id_stage_i/_0284_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1109_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0284_ ),
    .B1(\i_ibex/id_stage_i/_0281_ ),
    .A1(net730),
    .Y(\i_ibex/id_stage_i/_0285_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1110_  (.B(net1374),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0286_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0285_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1111_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net685),
    .Y(\i_ibex/alu_operand_b_ex [23]),
    .A2(\i_ibex/id_stage_i/_0286_ ),
    .A1(\i_ibex/id_stage_i/_0280_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1112_  (.Y(\i_ibex/id_stage_i/_0287_ ),
    .B(\i_ibex/rf_rdata_b [22]),
    .A_N(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1113_  (.A0(net730),
    .A1(net755),
    .S(net673),
    .X(\i_ibex/id_stage_i/_0288_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1114_  (.Y(\i_ibex/id_stage_i/_0289_ ),
    .A(net1332),
    .B(net731),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1115_  (.Y(\i_ibex/id_stage_i/_0290_ ),
    .B(net731),
    .A_N(net1332),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1116_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0289_ ),
    .A2(\i_ibex/id_stage_i/_0290_ ),
    .Y(\i_ibex/id_stage_i/_0291_ ),
    .B1(net1246));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1117_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1251),
    .C1(\i_ibex/id_stage_i/_0291_ ),
    .B1(\i_ibex/id_stage_i/_0288_ ),
    .A1(net731),
    .Y(\i_ibex/id_stage_i/_0292_ ),
    .A2(net1190));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1118_  (.B(net1374),
    .C(net1242),
    .Y(\i_ibex/id_stage_i/_0293_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0292_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/_1119_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net679),
    .Y(\i_ibex/alu_operand_b_ex [22]),
    .A2(\i_ibex/id_stage_i/_0293_ ),
    .A1(\i_ibex/id_stage_i/_0287_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1120_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0294_ ),
    .A(\i_ibex/instr_fetch_err ),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/_1121_  (.B(net694),
    .C(\i_ibex/id_stage_i/_0294_ ),
    .A(net704),
    .Y(\i_ibex/id_stage_i/_0295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/_1122_  (.A(\i_ibex/id_stage_i/id_fsm_q ),
    .B(\i_ibex/id_stage_i/_0295_ ),
    .Y(\i_ibex/id_stage_i/_0296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/_1123_  (.B(\i_ibex/id_stage_i/jump_set_dec ),
    .C(\i_ibex/id_stage_i/_0296_ ),
    .A(\i_ibex/id_stage_i/jump_in_dec ),
    .Y(\i_ibex/id_stage_i/_0297_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/_1124_  (.A(\i_ibex/id_stage_i/branch_jump_set_done_q ),
    .B(\i_ibex/id_stage_i/branch_set_raw ),
    .Y(\i_ibex/id_stage_i/_0298_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1125_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0297_ ),
    .A2(\i_ibex/id_stage_i/_0298_ ),
    .Y(\i_ibex/id_stage_i/branch_jump_set_done_d ),
    .B1(\i_ibex/instr_valid_clear ));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1126_  (.A(\i_ibex/id_stage_i/branch_set_raw ),
    .B(\i_ibex/id_stage_i/jump_set_$_AND__Y_B ),
    .X(\i_ibex/id_stage_i/branch_set ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1127_  (.A(\i_ibex/id_stage_i/branch_in_dec ),
    .B(\i_ibex/id_stage_i/_0296_ ),
    .X(\i_ibex/perf_branch ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1128_  (.A(\i_ibex/branch_decision ),
    .B(\i_ibex/perf_branch ),
    .X(\i_ibex/id_stage_i/branch_set_raw_d ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1129_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0299_ ),
    .A(\i_ibex/id_stage_i/flush_id ),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/_1130_  (.X(\i_ibex/id_stage_i/_0300_ ),
    .A(net706),
    .B(net694),
    .C(\i_ibex/id_stage_i/_0294_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1131_  (.Y(\i_ibex/id_stage_i/_0301_ ),
    .B(\i_ibex/lsu_resp_valid ),
    .A_N(\i_ibex/id_stage_i/instr_first_cycle_id_o_$_AND__Y_B ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/_1132_  (.B(net704),
    .C(\i_ibex/id_stage_i/_0301_ ),
    .A(\i_ibex/id_stage_i/lsu_req_dec ),
    .Y(\i_ibex/id_stage_i/_0302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1133_  (.B1(\i_ibex/id_stage_i/branch_in_dec ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0303_ ),
    .VSS(VSS),
    .A1(\i_ibex/branch_decision ),
    .A2(\i_ibex/id_stage_i/id_fsm_q ));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1134_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0304_ ),
    .A(\i_ibex/id_stage_i/id_fsm_q ),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/_1135_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/_0305_ ),
    .B(net369),
    .A(net370));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/_1136_  (.Y(\i_ibex/id_stage_i/_0306_ ),
    .B(\i_ibex/ex_valid ),
    .A_N(\i_ibex/id_stage_i/id_fsm_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/_1137_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/id_stage_i/_0306_ ),
    .C1(\i_ibex/id_stage_i/jump_in_dec ),
    .B1(\i_ibex/id_stage_i/_0305_ ),
    .A1(net371),
    .Y(\i_ibex/id_stage_i/_0307_ ),
    .A2(\i_ibex/id_stage_i/_0304_ ));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1138_  (.A0(\i_ibex/ex_valid ),
    .A1(\i_ibex/lsu_resp_valid ),
    .S(\i_ibex/id_stage_i/lsu_req_dec ),
    .X(\i_ibex/id_stage_i/_0308_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1139_  (.A(\i_ibex/id_stage_i/id_fsm_q ),
    .B(\i_ibex/id_stage_i/_0308_ ),
    .X(\i_ibex/id_stage_i/_0309_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/id_stage_i/_1140_  (.A2(\i_ibex/id_stage_i/_0307_ ),
    .A1(\i_ibex/id_stage_i/_0303_ ),
    .B1(\i_ibex/id_stage_i/_0309_ ),
    .X(\i_ibex/id_stage_i/_0310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/id_stage_i/_1141_  (.A(\i_ibex/id_stage_i/_0299_ ),
    .B(\i_ibex/id_stage_i/_0300_ ),
    .C(\i_ibex/id_stage_i/_0302_ ),
    .D(\i_ibex/id_stage_i/_0310_ ),
    .X(\i_ibex/instr_id_done ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/id_stage_i/_1142_  (.A(net618),
    .B(\i_ibex/instr_id_done ),
    .X(\i_ibex/csr_op_en ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1143_  (.B(net750),
    .C(net745),
    .Y(\i_ibex/id_stage_i/_0311_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net747));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1144_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0312_ ),
    .A(net755),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/_1145_  (.B(\i_ibex/csr_op [1]),
    .C(\i_ibex/id_stage_i/_0312_ ),
    .A(\i_ibex/csr_op [0]),
    .Y(\i_ibex/id_stage_i/_0313_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net753));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/_1146_  (.Y(\i_ibex/id_stage_i/_0314_ ),
    .A(\i_ibex/csr_op [0]),
    .B(\i_ibex/csr_op [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/_1147_  (.A(net745),
    .B(net750),
    .C(net753),
    .Y(\i_ibex/id_stage_i/_0315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/_1148_  (.A(net757),
    .B(net761),
    .C(net747),
    .D(net755),
    .X(\i_ibex/id_stage_i/_0316_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1149_  (.B(\i_ibex/id_stage_i/_0315_ ),
    .C(\i_ibex/id_stage_i/_0316_ ),
    .Y(\i_ibex/id_stage_i/_0317_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/_0314_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1150_  (.B1(\i_ibex/id_stage_i/_0317_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0318_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/_0311_ ),
    .A2(\i_ibex/id_stage_i/_0313_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1151_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0319_ ),
    .A(net734),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/_1152_  (.B(net744),
    .C(net741),
    .Y(\i_ibex/id_stage_i/_0320_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net731));
 sg13g2_nor3_1 \i_ibex/id_stage_i/_1153_  (.A(\i_ibex/id_stage_i/_0319_ ),
    .B(net754),
    .C(\i_ibex/id_stage_i/_0320_ ),
    .Y(\i_ibex/id_stage_i/_0321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/_1154_  (.A(net757),
    .B(net761),
    .C(net747),
    .D(net754),
    .Y(\i_ibex/id_stage_i/_0322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1155_  (.Y(\i_ibex/id_stage_i/_0323_ ),
    .A(\i_ibex/id_stage_i/_0315_ ),
    .B(\i_ibex/id_stage_i/_0322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/id_stage_i/_1156_  (.A(net734),
    .B(\i_ibex/id_stage_i/_0314_ ),
    .C(\i_ibex/id_stage_i/_0320_ ),
    .X(\i_ibex/id_stage_i/_0324_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/_1157_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/_0311_ ),
    .A2(\i_ibex/id_stage_i/_0323_ ),
    .Y(\i_ibex/id_stage_i/_0325_ ),
    .B1(\i_ibex/id_stage_i/_0324_ ));
 sg13g2_a21o_2 \i_ibex/id_stage_i/_1158_  (.A2(\i_ibex/id_stage_i/_0321_ ),
    .A1(\i_ibex/id_stage_i/_0318_ ),
    .B1(\i_ibex/id_stage_i/_0325_ ),
    .X(\i_ibex/id_stage_i/_0326_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/_1159_  (.X(\i_ibex/id_stage_i/csr_pipe_flush ),
    .A(net618),
    .B(\i_ibex/instr_id_done ),
    .C(\i_ibex/id_stage_i/_0326_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1160_  (.A(net372),
    .B(\i_ibex/id_stage_i/_0300_ ),
    .X(\i_ibex/div_en_ex ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/_1161_  (.Y(\i_ibex/id_stage_i/_0327_ ),
    .A(\i_ibex/id_stage_i/_0300_ ),
    .B(\i_ibex/id_stage_i/_0308_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/_1162_  (.A(net373),
    .B(net374),
    .Y(\i_ibex/id_stage_i/_0328_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1163_  (.A(\i_ibex/branch_decision ),
    .B(\i_ibex/id_stage_i/branch_in_dec ),
    .X(\i_ibex/id_stage_i/_0329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/_1164_  (.A(\i_ibex/id_stage_i/jump_in_dec ),
    .B(net375),
    .C(\i_ibex/id_stage_i/lsu_req_dec ),
    .D(\i_ibex/id_stage_i/_0329_ ),
    .Y(\i_ibex/id_stage_i/_0330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1165_  (.B1(\i_ibex/id_stage_i/_0330_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0331_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_valid ),
    .A2(\i_ibex/id_stage_i/_0328_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/_1166_  (.Y(\i_ibex/id_stage_i/_0332_ ),
    .B1(\i_ibex/id_stage_i/_0331_ ),
    .B2(\i_ibex/id_stage_i/_0296_ ),
    .A2(\i_ibex/id_stage_i/_0327_ ),
    .A1(\i_ibex/id_stage_i/id_fsm_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1167_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0000_ ),
    .A(\i_ibex/id_stage_i/_0332_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1168_  (.B1(net704),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0333_ ),
    .VSS(VSS),
    .A1(\i_ibex/illegal_csr_insn_id ),
    .A2(\i_ibex/id_stage_i/illegal_insn_dec ));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1169_  (.VDD(VDD),
    .Y(\i_ibex/illegal_insn_id ),
    .A(\i_ibex/id_stage_i/_0333_ ),
    .VSS(VSS));
 sg13g2_buf_2 fanout633 (.A(net634),
    .X(net633),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout632 (.A(net634),
    .X(net632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1172_  (.A0(\i_ibex/imd_val_q_ex [0]),
    .A1(net257),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1173_  (.A0(\i_ibex/imd_val_q_ex [10]),
    .A1(net258),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1174_  (.A0(\i_ibex/imd_val_q_ex [11]),
    .A1(net259),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1175_  (.A0(\i_ibex/imd_val_q_ex [12]),
    .A1(net260),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1176_  (.A0(\i_ibex/imd_val_q_ex [13]),
    .A1(net261),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1177_  (.A0(\i_ibex/imd_val_q_ex [14]),
    .A1(net262),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1178_  (.A0(\i_ibex/imd_val_q_ex [15]),
    .A1(net263),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1179_  (.A0(\i_ibex/imd_val_q_ex [16]),
    .A1(net264),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1180_  (.A0(\i_ibex/imd_val_q_ex [17]),
    .A1(net265),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1181_  (.A0(\i_ibex/imd_val_q_ex [18]),
    .A1(net266),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout631 (.A(net634),
    .X(net631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1183_  (.A0(\i_ibex/imd_val_q_ex [19]),
    .A1(net267),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1184_  (.A0(\i_ibex/imd_val_q_ex [1]),
    .A1(net268),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1185_  (.A0(\i_ibex/imd_val_q_ex [20]),
    .A1(net269),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1186_  (.A0(\i_ibex/imd_val_q_ex [21]),
    .A1(net270),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1187_  (.A0(\i_ibex/imd_val_q_ex [22]),
    .A1(net271),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1188_  (.A0(\i_ibex/imd_val_q_ex [23]),
    .A1(net272),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1189_  (.A0(\i_ibex/imd_val_q_ex [24]),
    .A1(net273),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1190_  (.A0(\i_ibex/imd_val_q_ex [25]),
    .A1(net274),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1191_  (.A0(\i_ibex/imd_val_q_ex [26]),
    .A1(net275),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1192_  (.A0(\i_ibex/imd_val_q_ex [27]),
    .A1(net276),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout630 (.A(\i_ibex/pc_mux_id [2]),
    .X(net630),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1194_  (.A0(\i_ibex/imd_val_q_ex [28]),
    .A1(net277),
    .S(net1512),
    .X(\i_ibex/id_stage_i/_0021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1195_  (.A0(\i_ibex/imd_val_q_ex [29]),
    .A1(net278),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1196_  (.A0(\i_ibex/imd_val_q_ex [2]),
    .A1(net279),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1197_  (.A0(\i_ibex/imd_val_q_ex [30]),
    .A1(net280),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1198_  (.A0(\i_ibex/imd_val_q_ex [31]),
    .A1(net281),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1199_  (.A0(\i_ibex/imd_val_q_ex [32]),
    .A1(net250),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1200_  (.A0(\i_ibex/imd_val_q_ex [33]),
    .A1(net251),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout629 (.A(\i_ibex/pc_mux_id [2]),
    .X(net629),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout628 (.A(\i_ibex/pc_mux_id [2]),
    .X(net628),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1203_  (.A0(\i_ibex/imd_val_q_ex [34]),
    .A1(net283),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1204_  (.A0(\i_ibex/imd_val_q_ex [35]),
    .A1(net284),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1205_  (.A0(\i_ibex/imd_val_q_ex [36]),
    .A1(net285),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1206_  (.A0(\i_ibex/imd_val_q_ex [37]),
    .A1(net286),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1207_  (.A0(\i_ibex/imd_val_q_ex [38]),
    .A1(net287),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1208_  (.A0(\i_ibex/imd_val_q_ex [39]),
    .A1(net288),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1209_  (.A0(\i_ibex/imd_val_q_ex [3]),
    .A1(net289),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1210_  (.A0(\i_ibex/imd_val_q_ex [40]),
    .A1(net290),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1211_  (.A0(\i_ibex/imd_val_q_ex [41]),
    .A1(net291),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1212_  (.A0(\i_ibex/imd_val_q_ex [42]),
    .A1(net292),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1213_  (.A0(\i_ibex/imd_val_q_ex [43]),
    .A1(net293),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(\i_ibex/pc_mux_id [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1215_  (.A0(\i_ibex/imd_val_q_ex [44]),
    .A1(net294),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1216_  (.A0(\i_ibex/imd_val_q_ex [45]),
    .A1(net295),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1217_  (.A0(\i_ibex/imd_val_q_ex [46]),
    .A1(net296),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1218_  (.A0(\i_ibex/imd_val_q_ex [47]),
    .A1(net297),
    .S(net1507),
    .X(\i_ibex/id_stage_i/_0042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1219_  (.A0(\i_ibex/imd_val_q_ex [48]),
    .A1(net298),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1220_  (.A0(\i_ibex/imd_val_q_ex [49]),
    .A1(net299),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1221_  (.A0(\i_ibex/imd_val_q_ex [4]),
    .A1(net300),
    .S(net1512),
    .X(\i_ibex/id_stage_i/_0045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1222_  (.A0(\i_ibex/imd_val_q_ex [50]),
    .A1(net301),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1223_  (.A0(\i_ibex/imd_val_q_ex [51]),
    .A1(net302),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1224_  (.A0(\i_ibex/imd_val_q_ex [52]),
    .A1(net303),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1225_  (.A0(\i_ibex/imd_val_q_ex [53]),
    .A1(net304),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1227_  (.A0(\i_ibex/imd_val_q_ex [54]),
    .A1(net305),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1228_  (.A0(\i_ibex/imd_val_q_ex [55]),
    .A1(net306),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1229_  (.A0(\i_ibex/imd_val_q_ex [56]),
    .A1(net307),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1230_  (.A0(\i_ibex/imd_val_q_ex [57]),
    .A1(net308),
    .S(net1507),
    .X(\i_ibex/id_stage_i/_0053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1231_  (.A0(\i_ibex/imd_val_q_ex [58]),
    .A1(net309),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1232_  (.A0(\i_ibex/imd_val_q_ex [59]),
    .A1(net310),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1233_  (.A0(\i_ibex/imd_val_q_ex [5]),
    .A1(net311),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1234_  (.A0(\i_ibex/imd_val_q_ex [60]),
    .A1(net312),
    .S(net1507),
    .X(\i_ibex/id_stage_i/_0057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1235_  (.A0(\i_ibex/imd_val_q_ex [61]),
    .A1(net313),
    .S(net1505),
    .X(\i_ibex/id_stage_i/_0058_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1236_  (.A0(\i_ibex/imd_val_q_ex [62]),
    .A1(net314),
    .S(net1506),
    .X(\i_ibex/id_stage_i/_0059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1237_  (.A0(\i_ibex/imd_val_q_ex [63]),
    .A1(net315),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0060_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1238_  (.A0(\i_ibex/imd_val_q_ex [64]),
    .A1(net316),
    .S(net1504),
    .X(\i_ibex/id_stage_i/_0061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1239_  (.A0(\i_ibex/imd_val_q_ex [65]),
    .A1(net317),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1240_  (.A0(\i_ibex/imd_val_q_ex [66]),
    .A1(net252),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1241_  (.A0(\i_ibex/imd_val_q_ex [67]),
    .A1(net253),
    .S(net1503),
    .X(\i_ibex/id_stage_i/_0064_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1242_  (.A0(\i_ibex/imd_val_q_ex [6]),
    .A1(net318),
    .S(net1509),
    .X(\i_ibex/id_stage_i/_0065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1243_  (.A0(\i_ibex/imd_val_q_ex [7]),
    .A1(net319),
    .S(net1510),
    .X(\i_ibex/id_stage_i/_0066_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1244_  (.A0(\i_ibex/imd_val_q_ex [8]),
    .A1(net320),
    .S(net1511),
    .X(\i_ibex/id_stage_i/_0067_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1245_  (.A0(\i_ibex/imd_val_q_ex [9]),
    .A1(net321),
    .S(net1508),
    .X(\i_ibex/id_stage_i/_0068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1246_  (.A(net706),
    .B(\i_ibex/id_stage_i/instr_first_cycle_id_o_$_AND__Y_B ),
    .X(\i_ibex/instr_first_cycle_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/_1247_  (.A(net784),
    .B_N(\i_ibex/id_stage_i/dret_insn_dec ),
    .Y(\i_ibex/id_stage_i/_0342_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/_1248_  (.A(\i_ibex/illegal_csr_insn_id ),
    .B(\i_ibex/id_stage_i/illegal_insn_dec ),
    .C(\i_ibex/instr_fetch_err ),
    .Y(\i_ibex/id_stage_i/_0343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1249_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0344_ ),
    .A(\i_ibex/id_stage_i/_0343_ ),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/_1250_  (.A(\i_ibex/id_stage_i/ebrk_insn ),
    .B(\i_ibex/id_stage_i/ecall_insn_dec ),
    .C(\i_ibex/id_stage_i/_0342_ ),
    .D(\i_ibex/id_stage_i/_0344_ ),
    .Y(\i_ibex/instr_perf_count_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1251_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0345_ ),
    .A(\i_ibex/id_stage_i/jump_set_$_AND__Y_B ),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/_1252_  (.A(\i_ibex/id_stage_i/_0345_ ),
    .B(\i_ibex/id_stage_i/_0297_ ),
    .Y(\i_ibex/id_stage_i/jump_set ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/_1253_  (.X(\i_ibex/lsu_req ),
    .A(\i_ibex/id_stage_i/lsu_req_dec ),
    .B(\i_ibex/id_stage_i/_0300_ ),
    .C(net696),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/_1254_  (.A(net376),
    .B(\i_ibex/id_stage_i/_0300_ ),
    .X(\i_ibex/mult_en_ex ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1255_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0346_ ),
    .A(\i_ibex/id_stage_i/lsu_req_dec ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1256_  (.B1(\i_ibex/ex_valid ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0347_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/_0346_ ),
    .A2(\i_ibex/id_stage_i/_0304_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/_1257_  (.B(\i_ibex/id_stage_i/id_fsm_q ),
    .C(\i_ibex/lsu_resp_valid ),
    .A(\i_ibex/id_stage_i/lsu_req_dec ),
    .Y(\i_ibex/id_stage_i/_0348_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_1258_  (.X(\i_ibex/perf_div_wait ),
    .A(\i_ibex/div_en_ex ),
    .B(\i_ibex/id_stage_i/_0347_ ),
    .C(\i_ibex/id_stage_i/_0348_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/_1259_  (.A(\i_ibex/id_stage_i/_0346_ ),
    .B(\i_ibex/lsu_resp_valid ),
    .C(\i_ibex/id_stage_i/_0295_ ),
    .Y(\i_ibex/perf_dside_wait ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_1260_  (.X(\i_ibex/rf_ren_a ),
    .A(net706),
    .B(\i_ibex/id_stage_i/rf_ren_a_dec ),
    .C(\i_ibex/id_stage_i/_0343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_1261_  (.X(\i_ibex/rf_ren_b ),
    .A(net706),
    .B(\i_ibex/id_stage_i/rf_ren_b_dec ),
    .C(\i_ibex/id_stage_i/_0343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout625 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_005_ ),
    .X(net625),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout624 (.A(\i_ibex/csr_restore_mret_id ),
    .X(net624),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1264_  (.A0(\i_ibex/result_ex [31]),
    .A1(\i_ibex/csr_rdata [31]),
    .S(net1364),
    .X(\i_ibex/rf_wdata_id [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1265_  (.A0(\i_ibex/result_ex [30]),
    .A1(\i_ibex/csr_rdata [30]),
    .S(net1364),
    .X(\i_ibex/rf_wdata_id [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1266_  (.A0(\i_ibex/result_ex [21]),
    .A1(\i_ibex/csr_rdata [21]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1267_  (.A0(\i_ibex/result_ex [20]),
    .A1(\i_ibex/csr_rdata [20]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1268_  (.A0(\i_ibex/result_ex [19]),
    .A1(\i_ibex/csr_rdata [19]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1269_  (.A0(\i_ibex/result_ex [18]),
    .A1(\i_ibex/csr_rdata [18]),
    .S(net1364),
    .X(\i_ibex/rf_wdata_id [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1270_  (.A0(\i_ibex/result_ex [17]),
    .A1(\i_ibex/csr_rdata [17]),
    .S(net1364),
    .X(\i_ibex/rf_wdata_id [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1271_  (.A0(\i_ibex/result_ex [16]),
    .A1(\i_ibex/csr_rdata [16]),
    .S(net1365),
    .X(\i_ibex/rf_wdata_id [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1272_  (.A0(\i_ibex/result_ex [15]),
    .A1(\i_ibex/csr_rdata [15]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1273_  (.A0(\i_ibex/result_ex [14]),
    .A1(\i_ibex/csr_rdata [14]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout623 (.A(\i_ibex/pc_mux_id [0]),
    .X(net623),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1275_  (.A0(\i_ibex/result_ex [13]),
    .A1(\i_ibex/csr_rdata [13]),
    .S(net1361),
    .X(\i_ibex/rf_wdata_id [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1276_  (.A0(\i_ibex/result_ex [12]),
    .A1(\i_ibex/csr_rdata [12]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1277_  (.A0(\i_ibex/result_ex [29]),
    .A1(\i_ibex/csr_rdata [29]),
    .S(net1365),
    .X(\i_ibex/rf_wdata_id [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1278_  (.A0(\i_ibex/result_ex [11]),
    .A1(\i_ibex/csr_rdata [11]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1279_  (.A0(\i_ibex/result_ex [10]),
    .A1(\i_ibex/csr_rdata [10]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1280_  (.A0(\i_ibex/result_ex [9]),
    .A1(\i_ibex/csr_rdata [9]),
    .S(net1361),
    .X(\i_ibex/rf_wdata_id [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1281_  (.A0(\i_ibex/result_ex [8]),
    .A1(\i_ibex/csr_rdata [8]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1282_  (.A0(\i_ibex/result_ex [7]),
    .A1(\i_ibex/csr_rdata [7]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1283_  (.A0(\i_ibex/result_ex [6]),
    .A1(\i_ibex/csr_rdata [6]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1284_  (.A0(\i_ibex/result_ex [5]),
    .A1(\i_ibex/csr_rdata [5]),
    .S(net1360),
    .X(\i_ibex/rf_wdata_id [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout622 (.A(\i_ibex/alu_operator_ex [1]),
    .X(net622),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1286_  (.A0(\i_ibex/result_ex [4]),
    .A1(\i_ibex/csr_rdata [4]),
    .S(net1361),
    .X(\i_ibex/rf_wdata_id [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1287_  (.A0(\i_ibex/result_ex [3]),
    .A1(\i_ibex/csr_rdata [3]),
    .S(net1362),
    .X(\i_ibex/rf_wdata_id [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1288_  (.A0(\i_ibex/result_ex [2]),
    .A1(\i_ibex/csr_rdata [2]),
    .S(net1362),
    .X(\i_ibex/rf_wdata_id [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1289_  (.A0(\i_ibex/result_ex [28]),
    .A1(\i_ibex/csr_rdata [28]),
    .S(net1362),
    .X(\i_ibex/rf_wdata_id [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1290_  (.A0(\i_ibex/result_ex [1]),
    .A1(\i_ibex/csr_rdata [1]),
    .S(net1362),
    .X(\i_ibex/rf_wdata_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/_1291_  (.A0(\i_ibex/result_ex [0]),
    .A1(\i_ibex/csr_rdata [0]),
    .S(net1362),
    .X(\i_ibex/rf_wdata_id [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1292_  (.A0(\i_ibex/result_ex [27]),
    .A1(\i_ibex/csr_rdata [27]),
    .S(net1362),
    .X(\i_ibex/rf_wdata_id [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1293_  (.A0(\i_ibex/result_ex [26]),
    .A1(\i_ibex/csr_rdata [26]),
    .S(net1364),
    .X(\i_ibex/rf_wdata_id [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1294_  (.A0(\i_ibex/result_ex [25]),
    .A1(\i_ibex/csr_rdata [25]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1295_  (.A0(\i_ibex/result_ex [24]),
    .A1(\i_ibex/csr_rdata [24]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1296_  (.A0(\i_ibex/result_ex [23]),
    .A1(\i_ibex/csr_rdata [23]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/_1297_  (.A0(\i_ibex/result_ex [22]),
    .A1(\i_ibex/csr_rdata [22]),
    .S(net1363),
    .X(\i_ibex/rf_wdata_id [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/_1298_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0353_ ),
    .A(\i_ibex/id_stage_i/rf_we_dec ),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/_1299_  (.X(\i_ibex/id_stage_i/_0354_ ),
    .A(net377),
    .B(\i_ibex/id_stage_i/_0304_ ),
    .C(\i_ibex/id_stage_i/_0328_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1300_  (.B1(\i_ibex/id_stage_i/_0300_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/_0355_ ),
    .VSS(VSS),
    .A1(\i_ibex/ex_valid ),
    .A2(\i_ibex/id_stage_i/_0328_ ));
 sg13g2_nor4_1 \i_ibex/id_stage_i/_1301_  (.A(\i_ibex/id_stage_i/_0353_ ),
    .B(\i_ibex/illegal_csr_insn_id ),
    .C(\i_ibex/id_stage_i/_0354_ ),
    .D(\i_ibex/id_stage_i/_0355_ ),
    .Y(\i_ibex/rf_we_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/_1302_  (.B1(\i_ibex/id_stage_i/_0302_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/stall_id ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/_0295_ ),
    .A2(\i_ibex/id_stage_i/_0310_ ));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/branch_jump_set_done_q_reg  (.CLK(clknet_leaf_87_clk_i_regs),
    .RESET_B(net1576),
    .D(\i_ibex/id_stage_i/branch_jump_set_done_d ),
    .Q_N(\i_ibex/id_stage_i/jump_set_$_AND__Y_B ),
    .Q(\i_ibex/id_stage_i/branch_jump_set_done_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/branch_set_raw_reg  (.CLK(clknet_leaf_89_clk_i_regs),
    .RESET_B(net1577),
    .D(\i_ibex/id_stage_i/branch_set_raw_d ),
    .Q_N(\i_ibex/id_stage_i/_0627_ ),
    .Q(\i_ibex/id_stage_i/branch_set_raw ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 \i_ibex/id_stage_i/controller_i/_407_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_006_ ),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__B_Y_$_OR__Y_A ),
    .A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_408_  (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .B(net1487),
    .C(\i_ibex/id_stage_i/controller_i/_006_ ),
    .Y(\i_ibex/id_stage_i/controller_run ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout621 (.A(\i_ibex/alu_operator_ex [1]),
    .X(net621),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_410_  (.A(net706),
    .B(\i_ibex/instr_fetch_err ),
    .X(\i_ibex/id_stage_i/controller_i/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout620 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_084_ ),
    .X(net620),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(\i_ibex/csr_access ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_413_  (.A(\i_ibex/pc_id [28]),
    .B(\i_ibex/pc_id [27]),
    .X(\i_ibex/id_stage_i/controller_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_414_  (.Y(\i_ibex/id_stage_i/controller_i/_012_ ),
    .A(\i_ibex/instr_fetch_err_plus2 ),
    .B(\i_ibex/pc_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_415_  (.B(\i_ibex/pc_id [4]),
    .C(\i_ibex/pc_id [3]),
    .A(\i_ibex/pc_id [5]),
    .Y(\i_ibex/id_stage_i/controller_i/_013_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/pc_id [2]));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_416_  (.Y(\i_ibex/id_stage_i/controller_i/_014_ ),
    .A(\i_ibex/pc_id [7]),
    .B(\i_ibex/pc_id [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_417_  (.A(\i_ibex/id_stage_i/controller_i/_012_ ),
    .B(\i_ibex/id_stage_i/controller_i/_013_ ),
    .C(\i_ibex/id_stage_i/controller_i/_014_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/controller_i/_418_  (.A(\i_ibex/pc_id [11]),
    .B(\i_ibex/pc_id [10]),
    .C(\i_ibex/pc_id [9]),
    .D(\i_ibex/pc_id [8]),
    .X(\i_ibex/id_stage_i/controller_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/controller_i/_419_  (.X(\i_ibex/id_stage_i/controller_i/_017_ ),
    .A(\i_ibex/pc_id [13]),
    .B(\i_ibex/pc_id [12]),
    .C(\i_ibex/id_stage_i/controller_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/controller_i/_420_  (.A(\i_ibex/pc_id [17]),
    .B(\i_ibex/pc_id [16]),
    .C(\i_ibex/pc_id [15]),
    .D(\i_ibex/pc_id [14]),
    .X(\i_ibex/id_stage_i/controller_i/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/controller_i/_421_  (.X(\i_ibex/id_stage_i/controller_i/_019_ ),
    .A(\i_ibex/id_stage_i/controller_i/_015_ ),
    .B(\i_ibex/id_stage_i/controller_i/_017_ ),
    .C(\i_ibex/id_stage_i/controller_i/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout618 (.A(net619),
    .X(net618),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_423_  (.B(\i_ibex/pc_id [19]),
    .C(\i_ibex/pc_id [18]),
    .A(\i_ibex/pc_id [20]),
    .Y(\i_ibex/id_stage_i/controller_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_424_  (.B(\i_ibex/pc_id [22]),
    .C(\i_ibex/pc_id [21]),
    .A(\i_ibex/pc_id [23]),
    .Y(\i_ibex/id_stage_i/controller_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_425_  (.A(\i_ibex/id_stage_i/controller_i/_021_ ),
    .B(\i_ibex/id_stage_i/controller_i/_022_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_426_  (.A(\i_ibex/pc_id [24]),
    .B(\i_ibex/id_stage_i/controller_i/_023_ ),
    .X(\i_ibex/id_stage_i/controller_i/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/id_stage_i/controller_i/_427_  (.A(\i_ibex/pc_id [26]),
    .B(\i_ibex/pc_id [25]),
    .C(\i_ibex/id_stage_i/controller_i/_019_ ),
    .D(\i_ibex/id_stage_i/controller_i/_024_ ),
    .X(\i_ibex/id_stage_i/controller_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_428_  (.B(\i_ibex/pc_id [29]),
    .C(\i_ibex/id_stage_i/controller_i/_011_ ),
    .A(\i_ibex/pc_id [30]),
    .Y(\i_ibex/id_stage_i/controller_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_025_ ));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_429_  (.Y(\i_ibex/id_stage_i/controller_i/_027_ ),
    .A(\i_ibex/pc_id [31]),
    .B(\i_ibex/id_stage_i/controller_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_430_  (.Y(\i_ibex/id_stage_i/controller_i/_028_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout617 (.A(net618),
    .X(net617),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_432_  (.A(\i_ibex/id_stage_i/controller_i/store_err_q ),
    .B(\i_ibex/id_stage_i/controller_i/load_err_q ),
    .Y(\i_ibex/id_stage_i/controller_i/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/id_stage_i/controller_i/_433_  (.Y(\i_ibex/id_stage_i/controller_i/_031_ ),
    .A(net704),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_434_  (.A(\i_ibex/id_stage_i/ebrk_insn ),
    .B(\i_ibex/id_stage_i/ecall_insn_dec ),
    .C(\i_ibex/instr_fetch_err ),
    .Y(\i_ibex/id_stage_i/controller_i/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_435_  (.A(\i_ibex/id_stage_i/controller_i/_031_ ),
    .B(\i_ibex/id_stage_i/controller_i/_032_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_436_  (.A(\i_ibex/id_stage_i/controller_i/illegal_insn_q ),
    .B(\i_ibex/id_stage_i/controller_i/_030_ ),
    .C(\i_ibex/id_stage_i/controller_i/_033_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout616 (.A(net618),
    .X(net616),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/id_stage_i/controller_i/_438_  (.Y(\i_ibex/id_stage_i/controller_i/_036_ ),
    .A(net1485),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout615 (.A(\i_ibex/id_stage_i/controller_i/_034_ ),
    .X(net615),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_440_  (.A(\i_ibex/id_stage_i/controller_i/_036_ ),
    .B(net783),
    .C(net1455),
    .Y(\i_ibex/id_stage_i/controller_i/_038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_442_  (.Y(\i_ibex/id_stage_i/controller_i/_040_ ),
    .B1(net1395),
    .B2(net731),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout613 (.A(net615),
    .X(net613),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_444_  (.A(net1489),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .C(\i_ibex/id_stage_i/controller_i/_006_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_445_  (.A(\i_ibex/id_stage_i/controller_i/exc_req_q ),
    .B(\i_ibex/id_stage_i/controller_i/store_err_q ),
    .C(\i_ibex/id_stage_i/controller_i/load_err_q ),
    .Y(\i_ibex/id_stage_i/controller_i/_043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_446_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_044_ ),
    .A(\i_ibex/id_stage_i/controller_i/_043_ ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_447_  (.Y(\i_ibex/id_stage_i/controller_i/_045_ ),
    .A(\i_ibex/id_stage_i/controller_i/_042_ ),
    .B(\i_ibex/id_stage_i/controller_i/_044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout612 (.A(net615),
    .X(net612),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout611 (.A(net615),
    .X(net611),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_450_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1407),
    .Y(\i_ibex/csr_mtval [31]),
    .A2(\i_ibex/id_stage_i/controller_i/_040_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_028_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_451_  (.B(\i_ibex/id_stage_i/controller_i/_011_ ),
    .C(\i_ibex/id_stage_i/controller_i/_025_ ),
    .A(\i_ibex/pc_id [29]),
    .Y(\i_ibex/id_stage_i/controller_i/_048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_452_  (.Y(\i_ibex/id_stage_i/controller_i/_049_ ),
    .A(\i_ibex/pc_id [30]),
    .B(\i_ibex/id_stage_i/controller_i/_048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_453_  (.Y(\i_ibex/id_stage_i/controller_i/_050_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_454_  (.Y(\i_ibex/id_stage_i/controller_i/_051_ ),
    .B1(net1396),
    .B2(net734),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_455_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1407),
    .Y(\i_ibex/csr_mtval [30]),
    .A2(\i_ibex/id_stage_i/controller_i/_051_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_050_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/controller_i/_456_  (.A(\i_ibex/id_stage_i/controller_i/_021_ ),
    .B_N(\i_ibex/id_stage_i/controller_i/_019_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_457_  (.B(\i_ibex/id_stage_i/controller_i/_052_ ),
    .A(\i_ibex/pc_id [21]),
    .X(\i_ibex/id_stage_i/controller_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_458_  (.Y(\i_ibex/id_stage_i/controller_i/_054_ ),
    .A(net1454),
    .B(\i_ibex/id_stage_i/controller_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_459_  (.Y(\i_ibex/id_stage_i/controller_i/_055_ ),
    .B1(net1395),
    .B2(net757),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_460_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1407),
    .Y(\i_ibex/csr_mtval [21]),
    .A2(\i_ibex/id_stage_i/controller_i/_055_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_054_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_461_  (.B(\i_ibex/pc_id [18]),
    .C(\i_ibex/id_stage_i/controller_i/_019_ ),
    .A(\i_ibex/pc_id [19]),
    .Y(\i_ibex/id_stage_i/controller_i/_056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_462_  (.Y(\i_ibex/id_stage_i/controller_i/_057_ ),
    .A(\i_ibex/pc_id [20]),
    .B(\i_ibex/id_stage_i/controller_i/_056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_463_  (.Y(\i_ibex/id_stage_i/controller_i/_058_ ),
    .A(net1455),
    .B(\i_ibex/id_stage_i/controller_i/_057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout610 (.A(\i_ibex/csr_save_if ),
    .X(net610),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_465_  (.Y(\i_ibex/id_stage_i/controller_i/_060_ ),
    .B1(net1396),
    .B2(net761),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_466_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1408),
    .Y(\i_ibex/csr_mtval [20]),
    .A2(\i_ibex/id_stage_i/controller_i/_060_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_058_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_467_  (.Y(\i_ibex/id_stage_i/controller_i/_061_ ),
    .A(\i_ibex/pc_id [18]),
    .B(\i_ibex/id_stage_i/controller_i/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_468_  (.Y(\i_ibex/id_stage_i/controller_i/_062_ ),
    .A(\i_ibex/pc_id [19]),
    .B(\i_ibex/id_stage_i/controller_i/_061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_469_  (.Y(\i_ibex/id_stage_i/controller_i/_063_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_470_  (.Y(\i_ibex/id_stage_i/controller_i/_064_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_038_ ),
    .B2(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_471_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_063_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_064_ ),
    .Y(\i_ibex/csr_mtval [19]),
    .B1(net1408));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_472_  (.B(\i_ibex/id_stage_i/controller_i/_019_ ),
    .A(\i_ibex/pc_id [18]),
    .X(\i_ibex/id_stage_i/controller_i/_065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_473_  (.Y(\i_ibex/id_stage_i/controller_i/_066_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_474_  (.Y(\i_ibex/id_stage_i/controller_i/_067_ ),
    .B1(net1395),
    .B2(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_475_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_066_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_067_ ),
    .Y(\i_ibex/csr_mtval [18]),
    .B1(net1406));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_476_  (.A(\i_ibex/id_stage_i/controller_i/_015_ ),
    .B(\i_ibex/id_stage_i/controller_i/_017_ ),
    .X(\i_ibex/id_stage_i/controller_i/_068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_477_  (.B(\i_ibex/pc_id [15]),
    .C(\i_ibex/pc_id [14]),
    .A(\i_ibex/pc_id [16]),
    .Y(\i_ibex/id_stage_i/controller_i/_069_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_068_ ));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_478_  (.Y(\i_ibex/id_stage_i/controller_i/_070_ ),
    .A(\i_ibex/pc_id [17]),
    .B(\i_ibex/id_stage_i/controller_i/_069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_479_  (.Y(\i_ibex/id_stage_i/controller_i/_071_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_070_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_480_  (.Y(\i_ibex/id_stage_i/controller_i/_072_ ),
    .B1(net1396),
    .B2(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_481_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_071_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_072_ ),
    .Y(\i_ibex/csr_mtval [17]),
    .B1(net1407));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_482_  (.B(\i_ibex/pc_id [14]),
    .C(\i_ibex/id_stage_i/controller_i/_068_ ),
    .A(\i_ibex/pc_id [15]),
    .Y(\i_ibex/id_stage_i/controller_i/_073_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_483_  (.Y(\i_ibex/id_stage_i/controller_i/_074_ ),
    .A(\i_ibex/pc_id [16]),
    .B(\i_ibex/id_stage_i/controller_i/_073_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_484_  (.Y(\i_ibex/id_stage_i/controller_i/_075_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_485_  (.Y(\i_ibex/id_stage_i/controller_i/_076_ ),
    .B1(net1396),
    .B2(net766),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_486_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1407),
    .Y(\i_ibex/csr_mtval [16]),
    .A2(\i_ibex/id_stage_i/controller_i/_076_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_075_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_487_  (.Y(\i_ibex/id_stage_i/controller_i/_077_ ),
    .A(\i_ibex/pc_id [14]),
    .B(\i_ibex/id_stage_i/controller_i/_068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_488_  (.Y(\i_ibex/id_stage_i/controller_i/_078_ ),
    .A(\i_ibex/pc_id [15]),
    .B(\i_ibex/id_stage_i/controller_i/_077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_489_  (.Y(\i_ibex/id_stage_i/controller_i/_079_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/controller_i/_490_  (.A(\i_ibex/id_stage_i/controller_i/_036_ ),
    .B(net1455),
    .Y(\i_ibex/id_stage_i/controller_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(net610),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_492_  (.A0(net768),
    .A1(\i_ibex/instr_rdata_c_id [15]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_493_  (.Y(\i_ibex/id_stage_i/controller_i/_083_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_082_ ),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_494_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1407),
    .Y(\i_ibex/csr_mtval [15]),
    .A2(\i_ibex/id_stage_i/controller_i/_083_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_079_ ));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_495_  (.B(\i_ibex/id_stage_i/controller_i/_068_ ),
    .A(\i_ibex/pc_id [14]),
    .X(\i_ibex/id_stage_i/controller_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_496_  (.Y(\i_ibex/id_stage_i/controller_i/_085_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_497_  (.A0(net770),
    .A1(\i_ibex/instr_rdata_c_id [14]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_498_  (.Y(\i_ibex/id_stage_i/controller_i/_087_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_086_ ),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_499_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1404),
    .Y(\i_ibex/csr_mtval [14]),
    .A2(\i_ibex/id_stage_i/controller_i/_087_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_085_ ));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net610),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_501_  (.B(\i_ibex/id_stage_i/controller_i/_015_ ),
    .C(\i_ibex/id_stage_i/controller_i/_016_ ),
    .A(\i_ibex/pc_id [12]),
    .Y(\i_ibex/id_stage_i/controller_i/_089_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_502_  (.Y(\i_ibex/id_stage_i/controller_i/_090_ ),
    .A(\i_ibex/pc_id [13]),
    .B(\i_ibex/id_stage_i/controller_i/_089_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_503_  (.Y(\i_ibex/id_stage_i/controller_i/_091_ ),
    .A(net1452),
    .B(\i_ibex/id_stage_i/controller_i/_090_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_504_  (.A0(net774),
    .A1(\i_ibex/instr_rdata_c_id [13]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_505_  (.Y(\i_ibex/id_stage_i/controller_i/_093_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_080_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_092_ ),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(net610),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_507_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1405),
    .Y(\i_ibex/csr_mtval [13]),
    .A2(\i_ibex/id_stage_i/controller_i/_093_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_091_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_508_  (.Y(\i_ibex/id_stage_i/controller_i/_095_ ),
    .A(\i_ibex/id_stage_i/controller_i/_015_ ),
    .B(\i_ibex/id_stage_i/controller_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_509_  (.Y(\i_ibex/id_stage_i/controller_i/_096_ ),
    .A(\i_ibex/pc_id [12]),
    .B(\i_ibex/id_stage_i/controller_i/_095_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_510_  (.Y(\i_ibex/id_stage_i/controller_i/_097_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_096_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_511_  (.A0(net778),
    .A1(\i_ibex/instr_rdata_c_id [12]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_512_  (.Y(\i_ibex/id_stage_i/controller_i/_099_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_080_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_098_ ),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_513_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1405),
    .Y(\i_ibex/csr_mtval [12]),
    .A2(\i_ibex/id_stage_i/controller_i/_099_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_097_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_514_  (.Y(\i_ibex/id_stage_i/controller_i/_100_ ),
    .A(\i_ibex/id_stage_i/controller_i/_011_ ),
    .B(\i_ibex/id_stage_i/controller_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_515_  (.Y(\i_ibex/id_stage_i/controller_i/_101_ ),
    .A(\i_ibex/pc_id [29]),
    .B(\i_ibex/id_stage_i/controller_i/_100_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_516_  (.Y(\i_ibex/id_stage_i/controller_i/_102_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_517_  (.Y(\i_ibex/id_stage_i/controller_i/_103_ ),
    .B1(net1396),
    .B2(net742),
    .A2(net612),
    .A1(\i_ibex/lsu_addr_last [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_518_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1405),
    .Y(\i_ibex/csr_mtval [29]),
    .A2(\i_ibex/id_stage_i/controller_i/_103_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_102_ ));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_519_  (.B(\i_ibex/pc_id [9]),
    .C(\i_ibex/pc_id [8]),
    .A(\i_ibex/pc_id [10]),
    .Y(\i_ibex/id_stage_i/controller_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_015_ ));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_520_  (.Y(\i_ibex/id_stage_i/controller_i/_105_ ),
    .A(\i_ibex/pc_id [11]),
    .B(\i_ibex/id_stage_i/controller_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_521_  (.Y(\i_ibex/id_stage_i/controller_i/_106_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(net610),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_523_  (.A0(\i_ibex/id_stage_i/imm_s_type [4]),
    .A1(\i_ibex/instr_rdata_c_id [11]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_524_  (.Y(\i_ibex/id_stage_i/controller_i/_109_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_108_ ),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_525_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1404),
    .Y(\i_ibex/csr_mtval [11]),
    .A2(\i_ibex/id_stage_i/controller_i/_109_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_106_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_526_  (.B(\i_ibex/pc_id [8]),
    .C(\i_ibex/id_stage_i/controller_i/_015_ ),
    .A(\i_ibex/pc_id [9]),
    .Y(\i_ibex/id_stage_i/controller_i/_110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_527_  (.Y(\i_ibex/id_stage_i/controller_i/_111_ ),
    .A(\i_ibex/pc_id [10]),
    .B(\i_ibex/id_stage_i/controller_i/_110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_528_  (.Y(\i_ibex/id_stage_i/controller_i/_112_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_529_  (.A0(\i_ibex/id_stage_i/imm_s_type [3]),
    .A1(\i_ibex/instr_rdata_c_id [10]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_530_  (.Y(\i_ibex/id_stage_i/controller_i/_114_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_113_ ),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_531_  (.Y(\i_ibex/id_stage_i/controller_i/_115_ ),
    .A(net705),
    .B(\i_ibex/instr_fetch_err ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_532_  (.Y(\i_ibex/id_stage_i/controller_i/_116_ ),
    .A(\i_ibex/id_stage_i/controller_i/_036_ ),
    .B(\i_ibex/id_stage_i/controller_i/_115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/id_stage_i/controller_i/_533_  (.A(net1490),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .C(\i_ibex/id_stage_i/controller_i/_006_ ),
    .X(\i_ibex/id_stage_i/controller_i/_117_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout605 (.A(\i_ibex/ex_block_i/alu_i/_0621_ ),
    .X(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/controller_i/_535_  (.A(net1449),
    .B(\i_ibex/id_stage_i/controller_i/_043_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_536_  (.B1(\i_ibex/id_stage_i/controller_i/_119_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_120_ ),
    .VSS(VSS),
    .A1(net615),
    .A2(\i_ibex/id_stage_i/controller_i/_116_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_537_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/controller_i/_120_ ),
    .Y(\i_ibex/csr_mtval [10]),
    .A2(\i_ibex/id_stage_i/controller_i/_114_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_112_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_538_  (.Y(\i_ibex/id_stage_i/controller_i/_121_ ),
    .A(\i_ibex/pc_id [8]),
    .B(\i_ibex/id_stage_i/controller_i/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_539_  (.Y(\i_ibex/id_stage_i/controller_i/_122_ ),
    .A(\i_ibex/pc_id [9]),
    .B(\i_ibex/id_stage_i/controller_i/_121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_540_  (.Y(\i_ibex/id_stage_i/controller_i/_123_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_541_  (.A0(\i_ibex/id_stage_i/imm_s_type [2]),
    .A1(\i_ibex/instr_rdata_c_id [9]),
    .S(net782),
    .X(\i_ibex/id_stage_i/controller_i/_124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_542_  (.Y(\i_ibex/id_stage_i/controller_i/_125_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_124_ ),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_543_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1404),
    .Y(\i_ibex/csr_mtval [9]),
    .A2(\i_ibex/id_stage_i/controller_i/_125_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_123_ ));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_544_  (.B(\i_ibex/id_stage_i/controller_i/_015_ ),
    .A(\i_ibex/pc_id [8]),
    .X(\i_ibex/id_stage_i/controller_i/_126_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_545_  (.Y(\i_ibex/id_stage_i/controller_i/_127_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_126_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_546_  (.A0(\i_ibex/id_stage_i/imm_s_type [1]),
    .A1(\i_ibex/instr_rdata_c_id [8]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_547_  (.Y(\i_ibex/id_stage_i/controller_i/_129_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_128_ ),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_548_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/controller_i/_120_ ),
    .Y(\i_ibex/csr_mtval [8]),
    .A2(\i_ibex/id_stage_i/controller_i/_129_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_127_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_549_  (.A(\i_ibex/id_stage_i/controller_i/_012_ ),
    .B(\i_ibex/id_stage_i/controller_i/_013_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_550_  (.Y(\i_ibex/id_stage_i/controller_i/_131_ ),
    .A(\i_ibex/pc_id [6]),
    .B(\i_ibex/id_stage_i/controller_i/_130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_551_  (.B(\i_ibex/id_stage_i/controller_i/_131_ ),
    .A(\i_ibex/pc_id [7]),
    .X(\i_ibex/id_stage_i/controller_i/_132_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_552_  (.A0(\i_ibex/id_stage_i/imm_s_type [0]),
    .A1(\i_ibex/instr_rdata_c_id [7]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_553_  (.Y(\i_ibex/id_stage_i/controller_i/_134_ ),
    .B1(net1394),
    .B2(\i_ibex/id_stage_i/controller_i/_133_ ),
    .A2(net611),
    .A1(\i_ibex/lsu_addr_last [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_554_  (.B1(\i_ibex/id_stage_i/controller_i/_134_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_135_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_115_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_132_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_555_  (.A(\i_ibex/id_stage_i/controller_i/_119_ ),
    .B(\i_ibex/id_stage_i/controller_i/_135_ ),
    .X(\i_ibex/csr_mtval [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout604 (.A(net605),
    .X(net604),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_557_  (.Y(\i_ibex/id_stage_i/controller_i/_137_ ),
    .A(\i_ibex/pc_id [6]),
    .B(\i_ibex/id_stage_i/controller_i/_130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_558_  (.A0(net708),
    .A1(\i_ibex/instr_rdata_c_id [6]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_138_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_559_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1485),
    .A2(\i_ibex/id_stage_i/controller_i/_138_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_139_ ),
    .B1(net1451));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_560_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1451),
    .A2(\i_ibex/id_stage_i/controller_i/_137_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_140_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_139_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_561_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/lsu_addr_last [6]),
    .A2(net611),
    .Y(\i_ibex/id_stage_i/controller_i/_141_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_140_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_562_  (.A(net1404),
    .B(\i_ibex/id_stage_i/controller_i/_141_ ),
    .Y(\i_ibex/csr_mtval [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_563_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_142_ ),
    .A(\i_ibex/id_stage_i/controller_i/_012_ ),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_564_  (.B(\i_ibex/pc_id [3]),
    .C(\i_ibex/pc_id [2]),
    .A(\i_ibex/pc_id [4]),
    .Y(\i_ibex/id_stage_i/controller_i/_143_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_142_ ));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_565_  (.B(\i_ibex/id_stage_i/controller_i/_143_ ),
    .A(\i_ibex/pc_id [5]),
    .X(\i_ibex/id_stage_i/controller_i/_144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_566_  (.A0(net712),
    .A1(\i_ibex/instr_rdata_c_id [5]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_567_  (.B(\i_ibex/id_stage_i/controller_i/_115_ ),
    .C(\i_ibex/id_stage_i/controller_i/_145_ ),
    .A(net1485),
    .Y(\i_ibex/id_stage_i/controller_i/_146_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_568_  (.B1(\i_ibex/id_stage_i/controller_i/_146_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_147_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_115_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_144_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_569_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/lsu_addr_last [5]),
    .A2(net611),
    .Y(\i_ibex/id_stage_i/controller_i/_148_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_147_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_570_  (.A(\i_ibex/id_stage_i/controller_i/_120_ ),
    .B(\i_ibex/id_stage_i/controller_i/_148_ ),
    .Y(\i_ibex/csr_mtval [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_571_  (.B(\i_ibex/pc_id [2]),
    .C(\i_ibex/id_stage_i/controller_i/_142_ ),
    .A(\i_ibex/pc_id [3]),
    .Y(\i_ibex/id_stage_i/controller_i/_149_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_572_  (.B(\i_ibex/id_stage_i/controller_i/_149_ ),
    .A(\i_ibex/pc_id [4]),
    .X(\i_ibex/id_stage_i/controller_i/_150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_573_  (.A0(net715),
    .A1(\i_ibex/instr_rdata_c_id [4]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_151_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_574_  (.B(\i_ibex/id_stage_i/controller_i/_115_ ),
    .C(\i_ibex/id_stage_i/controller_i/_151_ ),
    .A(net1485),
    .Y(\i_ibex/id_stage_i/controller_i/_152_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_575_  (.B1(\i_ibex/id_stage_i/controller_i/_152_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_153_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_115_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_150_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_576_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/lsu_addr_last [4]),
    .A2(net611),
    .Y(\i_ibex/id_stage_i/controller_i/_154_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_153_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_577_  (.A(net1404),
    .B(\i_ibex/id_stage_i/controller_i/_154_ ),
    .Y(\i_ibex/csr_mtval [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_578_  (.Y(\i_ibex/id_stage_i/controller_i/_155_ ),
    .A(\i_ibex/lsu_addr_last [3]),
    .B(net615),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_579_  (.Y(\i_ibex/id_stage_i/controller_i/_156_ ),
    .A(\i_ibex/pc_id [2]),
    .B(\i_ibex/id_stage_i/controller_i/_142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_580_  (.Y(\i_ibex/id_stage_i/controller_i/_157_ ),
    .A(\i_ibex/pc_id [3]),
    .B(\i_ibex/id_stage_i/controller_i/_156_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_581_  (.A0(net719),
    .A1(\i_ibex/instr_rdata_c_id [3]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_582_  (.Y(\i_ibex/id_stage_i/controller_i/_159_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_158_ ),
    .B2(net1394),
    .A2(\i_ibex/id_stage_i/controller_i/_157_ ),
    .A1(net1451),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_583_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1404),
    .Y(\i_ibex/csr_mtval [3]),
    .A2(\i_ibex/id_stage_i/controller_i/_159_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_155_ ));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_584_  (.B(\i_ibex/id_stage_i/controller_i/_012_ ),
    .A(\i_ibex/pc_id [2]),
    .X(\i_ibex/id_stage_i/controller_i/_160_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_585_  (.A0(net738),
    .A1(\i_ibex/instr_rdata_c_id [2]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_586_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1485),
    .A2(\i_ibex/id_stage_i/controller_i/_161_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_162_ ),
    .B1(net1451));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_587_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1452),
    .A2(\i_ibex/id_stage_i/controller_i/_160_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_163_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_162_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_588_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/lsu_addr_last [2]),
    .A2(net611),
    .Y(\i_ibex/id_stage_i/controller_i/_164_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_163_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_589_  (.A(net1404),
    .B(\i_ibex/id_stage_i/controller_i/_164_ ),
    .Y(\i_ibex/csr_mtval [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_590_  (.Y(\i_ibex/id_stage_i/controller_i/_165_ ),
    .A(\i_ibex/pc_id [27]),
    .B(\i_ibex/id_stage_i/controller_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_591_  (.Y(\i_ibex/id_stage_i/controller_i/_166_ ),
    .A(\i_ibex/pc_id [28]),
    .B(\i_ibex/id_stage_i/controller_i/_165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_592_  (.Y(\i_ibex/id_stage_i/controller_i/_167_ ),
    .A(net1453),
    .B(\i_ibex/id_stage_i/controller_i/_166_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_593_  (.Y(\i_ibex/id_stage_i/controller_i/_168_ ),
    .B1(net1396),
    .B2(net744),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_594_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1407),
    .Y(\i_ibex/csr_mtval [28]),
    .A2(\i_ibex/id_stage_i/controller_i/_168_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_167_ ));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_595_  (.Y(\i_ibex/id_stage_i/controller_i/_169_ ),
    .A(\i_ibex/instr_fetch_err_plus2 ),
    .B(\i_ibex/pc_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/id_stage_i/controller_i/_596_  (.A0(\i_ibex/instr_rdata_id [1]),
    .A1(\i_ibex/instr_rdata_c_id [1]),
    .S(net781),
    .X(\i_ibex/id_stage_i/controller_i/_170_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_597_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1485),
    .A2(\i_ibex/id_stage_i/controller_i/_170_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_171_ ),
    .B1(net1451));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_598_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1451),
    .A2(\i_ibex/id_stage_i/controller_i/_169_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_172_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_171_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_599_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/lsu_addr_last [1]),
    .A2(net611),
    .Y(\i_ibex/id_stage_i/controller_i/_173_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_172_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_600_  (.A(\i_ibex/id_stage_i/controller_i/_120_ ),
    .B(\i_ibex/id_stage_i/controller_i/_173_ ),
    .Y(\i_ibex/csr_mtval [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/controller_i/_601_  (.A(net783),
    .B_N(\i_ibex/instr_rdata_id [0]),
    .Y(\i_ibex/id_stage_i/controller_i/_174_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_602_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/controller_i/_174_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_175_ ),
    .A2(\i_ibex/instr_rdata_c_id [0]),
    .A1(net783));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_603_  (.A(\i_ibex/id_stage_i/controller_i/_036_ ),
    .B(net1451),
    .C(\i_ibex/id_stage_i/controller_i/_175_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/controller_i/_604_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/pc_id [0]),
    .C1(\i_ibex/id_stage_i/controller_i/_176_ ),
    .B1(net1451),
    .A1(\i_ibex/lsu_addr_last [0]),
    .Y(\i_ibex/id_stage_i/controller_i/_177_ ),
    .A2(net611));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_605_  (.A(net1404),
    .B(\i_ibex/id_stage_i/controller_i/_177_ ),
    .Y(\i_ibex/csr_mtval [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/id_stage_i/controller_i/_606_  (.B(\i_ibex/id_stage_i/controller_i/_025_ ),
    .A(\i_ibex/pc_id [27]),
    .X(\i_ibex/id_stage_i/controller_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_607_  (.Y(\i_ibex/id_stage_i/controller_i/_179_ ),
    .A(net1450),
    .B(\i_ibex/id_stage_i/controller_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_608_  (.Y(\i_ibex/id_stage_i/controller_i/_180_ ),
    .B1(net1396),
    .B2(net746),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_609_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1405),
    .Y(\i_ibex/csr_mtval [27]),
    .A2(\i_ibex/id_stage_i/controller_i/_180_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_179_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_610_  (.B(\i_ibex/id_stage_i/controller_i/_019_ ),
    .C(\i_ibex/id_stage_i/controller_i/_024_ ),
    .A(\i_ibex/pc_id [25]),
    .Y(\i_ibex/id_stage_i/controller_i/_181_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_611_  (.Y(\i_ibex/id_stage_i/controller_i/_182_ ),
    .A(\i_ibex/pc_id [26]),
    .B(\i_ibex/id_stage_i/controller_i/_181_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_612_  (.Y(\i_ibex/id_stage_i/controller_i/_183_ ),
    .A(net1454),
    .B(\i_ibex/id_stage_i/controller_i/_182_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_613_  (.Y(\i_ibex/id_stage_i/controller_i/_184_ ),
    .B1(net1395),
    .B2(net748),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_614_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1406),
    .Y(\i_ibex/csr_mtval [26]),
    .A2(\i_ibex/id_stage_i/controller_i/_184_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_183_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_615_  (.Y(\i_ibex/id_stage_i/controller_i/_185_ ),
    .A(\i_ibex/id_stage_i/controller_i/_019_ ),
    .B(\i_ibex/id_stage_i/controller_i/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_616_  (.Y(\i_ibex/id_stage_i/controller_i/_186_ ),
    .A(\i_ibex/pc_id [25]),
    .B(\i_ibex/id_stage_i/controller_i/_185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_617_  (.Y(\i_ibex/id_stage_i/controller_i/_187_ ),
    .A(net1454),
    .B(\i_ibex/id_stage_i/controller_i/_186_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_618_  (.Y(\i_ibex/id_stage_i/controller_i/_188_ ),
    .B1(net1395),
    .B2(net752),
    .A2(net614),
    .A1(\i_ibex/lsu_addr_last [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_619_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1406),
    .Y(\i_ibex/csr_mtval [25]),
    .A2(\i_ibex/id_stage_i/controller_i/_188_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_187_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_620_  (.Y(\i_ibex/id_stage_i/controller_i/_189_ ),
    .A(\i_ibex/id_stage_i/controller_i/_023_ ),
    .B(\i_ibex/id_stage_i/controller_i/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_621_  (.Y(\i_ibex/id_stage_i/controller_i/_190_ ),
    .A(\i_ibex/pc_id [24]),
    .B(\i_ibex/id_stage_i/controller_i/_189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_622_  (.Y(\i_ibex/id_stage_i/controller_i/_191_ ),
    .A(net1454),
    .B(\i_ibex/id_stage_i/controller_i/_190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_623_  (.Y(\i_ibex/id_stage_i/controller_i/_192_ ),
    .B1(net1395),
    .B2(net753),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_624_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1406),
    .Y(\i_ibex/csr_mtval [24]),
    .A2(\i_ibex/id_stage_i/controller_i/_192_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_191_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_625_  (.B(\i_ibex/pc_id [21]),
    .C(\i_ibex/id_stage_i/controller_i/_052_ ),
    .A(\i_ibex/pc_id [22]),
    .Y(\i_ibex/id_stage_i/controller_i/_193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_626_  (.Y(\i_ibex/id_stage_i/controller_i/_194_ ),
    .A(\i_ibex/pc_id [23]),
    .B(\i_ibex/id_stage_i/controller_i/_193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_627_  (.Y(\i_ibex/id_stage_i/controller_i/_195_ ),
    .A(net1455),
    .B(\i_ibex/id_stage_i/controller_i/_194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_628_  (.Y(\i_ibex/id_stage_i/controller_i/_196_ ),
    .B1(net1395),
    .B2(net754),
    .A2(net613),
    .A1(\i_ibex/lsu_addr_last [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_629_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1406),
    .Y(\i_ibex/csr_mtval [23]),
    .A2(\i_ibex/id_stage_i/controller_i/_196_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_195_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_630_  (.Y(\i_ibex/id_stage_i/controller_i/_197_ ),
    .A(\i_ibex/pc_id [21]),
    .B(\i_ibex/id_stage_i/controller_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/id_stage_i/controller_i/_631_  (.Y(\i_ibex/id_stage_i/controller_i/_198_ ),
    .A(\i_ibex/pc_id [22]),
    .B(\i_ibex/id_stage_i/controller_i/_197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_632_  (.Y(\i_ibex/id_stage_i/controller_i/_199_ ),
    .A(net1455),
    .B(\i_ibex/id_stage_i/controller_i/_198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_633_  (.Y(\i_ibex/id_stage_i/controller_i/_200_ ),
    .B1(net1395),
    .B2(net755),
    .A2(net611),
    .A1(\i_ibex/lsu_addr_last [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_634_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1406),
    .Y(\i_ibex/csr_mtval [22]),
    .A2(\i_ibex/id_stage_i/controller_i/_200_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_199_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_635_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_201_ ),
    .A(\i_ibex/id_stage_i/dret_insn_dec ),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_636_  (.Y(\i_ibex/id_stage_i/controller_i/_202_ ),
    .A(net705),
    .B(\i_ibex/id_stage_i/controller_i/_043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/id_stage_i/controller_i/_637_  (.A(\i_ibex/id_stage_i/controller_i/_201_ ),
    .B(\i_ibex/id_stage_i/mret_insn_dec ),
    .C(net1449),
    .Y(\i_ibex/csr_restore_dret_id ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_202_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_638_  (.A(net1449),
    .B(\i_ibex/id_stage_i/controller_i/_202_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_639_  (.Y(\i_ibex/id_stage_i/controller_i/_204_ ),
    .A(\i_ibex/id_stage_i/mret_insn_dec ),
    .B(\i_ibex/id_stage_i/controller_i/_203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_640_  (.VDD(VDD),
    .Y(\i_ibex/csr_restore_mret_id ),
    .A(\i_ibex/id_stage_i/controller_i/_204_ ),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_641_  (.A(\i_ibex/id_stage_i/controller_i/_031_ ),
    .B(net1485),
    .C(\i_ibex/instr_fetch_err ),
    .Y(\i_ibex/id_stage_i/controller_i/_205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/controller_i/_642_  (.B(\i_ibex/id_stage_i/controller_i/_205_ ),
    .C(\i_ibex/id_stage_i/ebrk_insn ),
    .Y(\i_ibex/id_stage_i/controller_i/_206_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/ecall_insn_dec ));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_643_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_207_ ),
    .A(net784),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_644_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_208_ ),
    .A(net786),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/controller_i/_645_  (.A(net785),
    .B_N(\i_ibex/debug_ebreaku ),
    .Y(\i_ibex/id_stage_i/controller_i/_209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_646_  (.Y(\i_ibex/id_stage_i/controller_i/_210_ ),
    .A(\i_ibex/id_stage_i/controller_i/_208_ ),
    .B(\i_ibex/id_stage_i/controller_i/_209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_647_  (.B(net785),
    .C(net786),
    .A(\i_ibex/debug_ebreakm ),
    .Y(\i_ibex/id_stage_i/controller_i/_211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/controller_i/_648_  (.X(\i_ibex/id_stage_i/controller_i/_212_ ),
    .A(\i_ibex/id_stage_i/controller_i/_207_ ),
    .B(\i_ibex/id_stage_i/controller_i/_210_ ),
    .C(\i_ibex/id_stage_i/controller_i/_211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_649_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_213_ ),
    .B(\i_ibex/id_stage_i/controller_i/_212_ ),
    .A(\i_ibex/id_stage_i/controller_i/_206_ ));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_651_  (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .B(net1486),
    .C(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ),
    .Y(\i_ibex/id_stage_i/controller_i/_215_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(\i_ibex/ex_block_i/alu_i/_0621_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_653_  (.A(net1487),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .C(\i_ibex/id_stage_i/controller_i/_006_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_217_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_654_  (.Y(\i_ibex/id_stage_i/controller_i/_218_ ),
    .A(net1489),
    .B(net1487),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_655_  (.B1(\i_ibex/id_stage_i/controller_i/_218_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_219_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_215_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_217_ ));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(\i_ibex/ex_block_i/alu_i/_0621_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_657_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_221_ ),
    .A(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_658_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_222_ ),
    .A(\i_ibex/id_stage_i/controller_i/_215_ ),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/id_stage_i/controller_i/_659_  (.A(\i_ibex/priv_mode_id [1]),
    .B(\i_ibex/priv_mode_id [0]),
    .X(\i_ibex/id_stage_i/controller_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_660_  (.Y(\i_ibex/id_stage_i/controller_i/_224_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_223_ ),
    .B2(\i_ibex/debug_ebreakm ),
    .A2(\i_ibex/id_stage_i/controller_i/_209_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_208_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/id_stage_i/controller_i/_661_  (.A(\i_ibex/id_stage_i/controller_i/_221_ ),
    .B(net1487),
    .C(\i_ibex/id_stage_i/controller_i/_222_ ),
    .D(\i_ibex/id_stage_i/controller_i/_224_ ),
    .X(\i_ibex/id_stage_i/controller_i/_225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_662_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/irq_pending_o ),
    .A2(\i_ibex/csr_mstatus_mie ),
    .Y(\i_ibex/id_stage_i/controller_i/_226_ ),
    .B1(net37));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/controller_i/_663_  (.A(\i_ibex/id_stage_i/controller_i/_226_ ),
    .B_N(\i_ibex/id_stage_i/controller_i/handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .Y(\i_ibex/id_stage_i/controller_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/id_stage_i/controller_i/_664_  (.A(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .B(\i_ibex/id_stage_i/controller_i/_227_ ),
    .X(\i_ibex/id_stage_i/controller_i/_228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_665_  (.Y(\i_ibex/id_stage_i/controller_i/_229_ ),
    .A(\i_ibex/id_stage_i/controller_i/_217_ ),
    .B(\i_ibex/id_stage_i/controller_i/_228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_666_  (.B1(\i_ibex/id_stage_i/controller_i/_229_ ),
    .VDD(VDD),
    .Y(\i_ibex/csr_save_if ),
    .VSS(VSS),
    .A1(net1489),
    .A2(\i_ibex/id_stage_i/controller_i/_222_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_667_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_230_ ),
    .A(\i_ibex/csr_save_if ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_668_  (.Y(\i_ibex/id_stage_i/controller_i/_231_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_225_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_230_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_219_ ),
    .A1(net1448),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/id_stage_i/controller_i/_669_  (.A2(\i_ibex/id_stage_i/controller_i/_213_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_119_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_231_ ),
    .X(\i_ibex/csr_save_cause ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_670_  (.VDD(VDD),
    .Y(\i_ibex/csr_save_id ),
    .A(\i_ibex/id_stage_i/controller_i/_225_ ),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_671_  (.A(debug_req_i),
    .B(net38),
    .Y(\i_ibex/id_stage_i/controller_i/_232_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_672_  (.A(\i_ibex/irq_pending_o ),
    .B(net784),
    .C(\i_ibex/debug_single_step ),
    .Y(\i_ibex/id_stage_i/controller_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_673_  (.Y(\i_ibex/id_stage_i/controller_i/_234_ ),
    .A(\i_ibex/id_stage_i/controller_i/_232_ ),
    .B(\i_ibex/id_stage_i/controller_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_674_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_235_ ),
    .A(net1490),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_675_  (.Y(\i_ibex/id_stage_i/controller_i/_236_ ),
    .A(\i_ibex/id_stage_i/controller_i/_235_ ),
    .B(net1488),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_676_  (.B1(\i_ibex/id_stage_i/controller_i/_236_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_237_ ),
    .VSS(VSS),
    .A1(net1488),
    .A2(\i_ibex/id_stage_i/controller_i/_234_ ));
 sg13g2_nor3_2 \i_ibex/id_stage_i/controller_i/_677_  (.A(net1486),
    .B(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .C(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .Y(\i_ibex/id_stage_i/controller_i/_238_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_678_  (.Y(\i_ibex/ctrl_busy ),
    .A(\i_ibex/id_stage_i/controller_i/_237_ ),
    .B(\i_ibex/id_stage_i/controller_i/_238_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_679_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_239_ ),
    .B(net1738),
    .A(\i_ibex/trigger_match ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_680_  (.A(\i_ibex/id_stage_i/controller_i/do_single_step_q ),
    .B(\i_ibex/id_stage_i/controller_i/_239_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_240_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_681_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_241_ ),
    .A(\i_ibex/id_stage_i/stall_id ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_682_  (.Y(\i_ibex/id_stage_i/controller_i/_242_ ),
    .A(\i_ibex/id_stage_i/controller_i/_031_ ),
    .B(\i_ibex/id_stage_i/controller_i/_241_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_683_  (.A(\i_ibex/id_stage_i/controller_i/_221_ ),
    .B(\i_ibex/id_stage_i/controller_i/_240_ ),
    .C(\i_ibex/id_stage_i/controller_i/_242_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_243_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_684_  (.A(net705),
    .B(\i_ibex/id_stage_i/stall_id ),
    .Y(\i_ibex/id_stage_i/controller_i/_244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_685_  (.B1(net705),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_245_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/csr_pipe_flush ),
    .A2(\i_ibex/perf_wfi_wait ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_686_  (.Y(\i_ibex/id_stage_i/controller_i/_246_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_245_ ),
    .B2(net1490),
    .A2(\i_ibex/id_stage_i/controller_i/_244_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/controller_i/_687_  (.A(\i_ibex/id_stage_i/dret_insn_dec ),
    .B(\i_ibex/id_stage_i/mret_insn_dec ),
    .Y(\i_ibex/id_stage_i/controller_i/_247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_688_  (.A(\i_ibex/id_stage_i/controller_i/_031_ ),
    .B(\i_ibex/id_stage_i/controller_i/_247_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_248_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/controller_i/_689_  (.A(\i_ibex/lsu_store_err ),
    .B(\i_ibex/lsu_load_err ),
    .Y(\i_ibex/id_stage_i/controller_i/_249_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_690_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/csr_mstatus_tw ),
    .A2(\i_ibex/perf_wfi_wait ),
    .Y(\i_ibex/id_stage_i/controller_i/_250_ ),
    .B1(\i_ibex/id_stage_i/mret_insn_dec ));
 sg13g2_or3_1 \i_ibex/id_stage_i/controller_i/_691_  (.A(\i_ibex/id_stage_i/controller_i/_031_ ),
    .B(\i_ibex/id_stage_i/controller_i/_223_ ),
    .C(\i_ibex/id_stage_i/controller_i/_250_ ),
    .X(\i_ibex/id_stage_i/controller_i/_251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_692_  (.B(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .C(\i_ibex/id_stage_i/dret_insn_dec ),
    .A(net704),
    .Y(\i_ibex/id_stage_i/controller_i/_252_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/controller_i/_693_  (.A(\i_ibex/illegal_insn_id ),
    .B_N(\i_ibex/id_stage_i/controller_i/_252_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/controller_i/_694_  (.B(\i_ibex/id_stage_i/controller_i/_251_ ),
    .C(\i_ibex/id_stage_i/controller_i/_253_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/controller_i/_033_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_695_  (.Y(\i_ibex/id_stage_i/controller_i/_255_ ),
    .A(net1448),
    .B(\i_ibex/id_stage_i/controller_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_696_  (.B(\i_ibex/id_stage_i/controller_i/_249_ ),
    .C(\i_ibex/id_stage_i/controller_i/_255_ ),
    .A(net694),
    .Y(\i_ibex/id_stage_i/controller_i/_256_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/id_stage_i/controller_i/_697_  (.A(\i_ibex/id_stage_i/controller_i/_243_ ),
    .B(\i_ibex/id_stage_i/controller_i/_246_ ),
    .C(\i_ibex/id_stage_i/controller_i/_248_ ),
    .D(\i_ibex/id_stage_i/controller_i/_256_ ),
    .X(\i_ibex/id_stage_i/controller_i/_257_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_698_  (.B1(\i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_q ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_258_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_224_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_206_ ));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_699_  (.B(\i_ibex/perf_wfi_wait ),
    .C(\i_ibex/id_stage_i/controller_i/_043_ ),
    .A(net707),
    .Y(\i_ibex/id_stage_i/controller_i/_259_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_247_ ));
 sg13g2_and3_1 \i_ibex/id_stage_i/controller_i/_700_  (.X(\i_ibex/id_stage_i/controller_i/_260_ ),
    .A(\i_ibex/id_stage_i/controller_i/_042_ ),
    .B(\i_ibex/id_stage_i/controller_i/_258_ ),
    .C(\i_ibex/id_stage_i/controller_i/_259_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_701_  (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [2]),
    .B(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .Y(\i_ibex/id_stage_i/controller_i/_261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_702_  (.Y(\i_ibex/id_stage_i/controller_i/_262_ ),
    .A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_703_  (.Y(\i_ibex/id_stage_i/controller_i/_263_ ),
    .A(\i_ibex/id_stage_i/controller_i/_261_ ),
    .B(\i_ibex/id_stage_i/controller_i/_262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_704_  (.A(net1490),
    .B(\i_ibex/id_stage_i/controller_i/_263_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_705_  (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__B_Y_$_OR__Y_A ),
    .Y(\i_ibex/id_stage_i/controller_i/_265_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/controller_i/_706_  (.A(net1489),
    .B(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .Y(\i_ibex/id_stage_i/controller_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_707_  (.A(\i_ibex/id_stage_i/controller_i/_265_ ),
    .B(\i_ibex/id_stage_i/controller_i/_266_ ),
    .X(\i_ibex/id_stage_i/controller_i/_267_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_708_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_268_ ),
    .A(\i_ibex/id_stage_i/controller_i/_267_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/id_stage_i/controller_i/_709_  (.A0(\i_ibex/id_stage_i/controller_i/do_single_step_q ),
    .A1(\i_ibex/debug_single_step ),
    .S(net706),
    .X(\i_ibex/id_stage_i/controller_i/_269_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_710_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_270_ ),
    .B(\i_ibex/id_stage_i/controller_i/_269_ ),
    .A(\i_ibex/id_stage_i/controller_i/_239_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_711_  (.Y(\i_ibex/id_stage_i/controller_i/_271_ ),
    .A(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .B(\i_ibex/id_stage_i/controller_i/_270_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_712_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_272_ ),
    .A(\i_ibex/id_stage_i/controller_i/_271_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_713_  (.B1(\i_ibex/id_stage_i/controller_i/_219_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_273_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_268_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_272_ ));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_714_  (.A(\i_ibex/id_stage_i/controller_i/_260_ ),
    .B(\i_ibex/id_stage_i/controller_i/_264_ ),
    .C(\i_ibex/id_stage_i/controller_i/_273_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_715_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .A2(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ),
    .Y(\i_ibex/id_stage_i/controller_i/_275_ ),
    .B1(net1486));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_716_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_276_ ),
    .A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_717_  (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .Y(\i_ibex/id_stage_i/controller_i/_277_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_718_  (.A(\i_ibex/id_stage_i/controller_i/_276_ ),
    .B(\i_ibex/id_stage_i/controller_i/_277_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_719_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1490),
    .A2(net1487),
    .Y(\i_ibex/id_stage_i/controller_i/_279_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_278_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_720_  (.B1(\i_ibex/id_stage_i/controller_i/_279_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_280_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_265_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_275_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_721_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_257_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_274_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_281_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_280_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_722_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1486),
    .A2(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__B_Y_$_OR__Y_A ),
    .Y(\i_ibex/id_stage_i/controller_i/_282_ ),
    .B1(net1489));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_723_  (.A(net1486),
    .B(net1487),
    .Y(\i_ibex/id_stage_i/controller_i/_283_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_724_  (.B1(\i_ibex/id_stage_i/controller_i/_277_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_284_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_282_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_283_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_725_  (.B(net1448),
    .C(\i_ibex/id_stage_i/controller_i/_254_ ),
    .A(net694),
    .Y(\i_ibex/id_stage_i/controller_i/_285_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/id_stage_i/controller_i/_726_  (.A(\i_ibex/id_stage_i/csr_pipe_flush ),
    .B(\i_ibex/id_stage_i/dret_insn_dec ),
    .C(\i_ibex/id_stage_i/mret_insn_dec ),
    .Y(\i_ibex/id_stage_i/controller_i/_286_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/perf_wfi_wait ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_727_  (.Y(\i_ibex/id_stage_i/controller_i/_287_ ),
    .B(net704),
    .A_N(\i_ibex/id_stage_i/controller_i/_286_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_728_  (.Y(\i_ibex/id_stage_i/controller_i/_288_ ),
    .A(\i_ibex/id_stage_i/controller_i/_249_ ),
    .B(\i_ibex/id_stage_i/controller_i/_287_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_729_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/stall_id ),
    .Y(\i_ibex/id_stage_i/controller_i/_289_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_288_ ),
    .A1(net694));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_730_  (.A(\i_ibex/id_stage_i/controller_i/_235_ ),
    .B(\i_ibex/id_stage_i/controller_i/_242_ ),
    .C(\i_ibex/id_stage_i/controller_i/_249_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_290_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_731_  (.B1(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_291_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_227_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_270_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_732_  (.B(\i_ibex/id_stage_i/controller_i/_265_ ),
    .C(\i_ibex/id_stage_i/controller_i/_218_ ),
    .A(\i_ibex/id_stage_i/controller_i/_276_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_292_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/id_stage_i/controller_i/_733_  (.A(\i_ibex/id_stage_i/controller_i/_290_ ),
    .B(\i_ibex/id_stage_i/controller_i/_291_ ),
    .C(\i_ibex/id_stage_i/controller_i/_292_ ),
    .X(\i_ibex/id_stage_i/controller_i/_293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/id_stage_i/controller_i/_734_  (.A(\i_ibex/id_stage_i/controller_i/_284_ ),
    .B(\i_ibex/id_stage_i/controller_i/_285_ ),
    .C(\i_ibex/id_stage_i/controller_i/_289_ ),
    .D(\i_ibex/id_stage_i/controller_i/_293_ ),
    .X(\i_ibex/id_in_ready ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_735_  (.Y(\i_ibex/id_stage_i/controller_i/_294_ ),
    .A(\i_ibex/id_stage_i/controller_i/_267_ ),
    .B(\i_ibex/id_stage_i/controller_i/_291_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_736_  (.A(net1490),
    .B(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .C(net1784),
    .Y(\i_ibex/id_stage_i/controller_i/_295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_737_  (.A(net1488),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .C(\i_ibex/id_stage_i/controller_i/_234_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_738_  (.B1(\i_ibex/id_stage_i/controller_i/_261_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_297_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_295_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_296_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_739_  (.B1(\i_ibex/id_stage_i/controller_i/_297_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_298_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_in_ready ),
    .A2(\i_ibex/id_stage_i/controller_i/_294_ ));
 sg13g2_mux2_1 \i_ibex/id_stage_i/controller_i/_740_  (.A0(\i_ibex/id_stage_i/controller_i/_281_ ),
    .A1(net1490),
    .S(\i_ibex/id_stage_i/controller_i/_298_ ),
    .X(\i_ibex/id_stage_i/controller_i/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_741_  (.B(\i_ibex/id_stage_i/controller_i/_203_ ),
    .C(\i_ibex/id_stage_i/controller_i/_258_ ),
    .A(\i_ibex/perf_wfi_wait ),
    .Y(\i_ibex/id_stage_i/controller_i/_299_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_247_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_742_  (.A(\i_ibex/id_stage_i/controller_i/_268_ ),
    .B(\i_ibex/id_stage_i/controller_i/_272_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_743_  (.A(net1489),
    .B(net1486),
    .Y(\i_ibex/id_stage_i/controller_i/_301_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_744_  (.Y(\i_ibex/id_stage_i/controller_i/_302_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_301_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_277_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_300_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_228_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/controller_i/_745_  (.A2(\i_ibex/id_stage_i/controller_i/_302_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_299_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_280_ ),
    .X(\i_ibex/id_stage_i/controller_i/_303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_746_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_251_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_253_ ),
    .Y(\i_ibex/id_stage_i/controller_i/illegal_insn_d ),
    .B1(\i_ibex/id_stage_i/controller_i/_042_ ));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/controller_i/_747_  (.B(\i_ibex/id_stage_i/controller_i/_249_ ),
    .C(\i_ibex/id_stage_i/controller_i/_243_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_304_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/controller_i/illegal_insn_d ));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_748_  (.A(net694),
    .B(\i_ibex/id_stage_i/controller_i/_304_ ),
    .X(\i_ibex/id_stage_i/controller_i/_305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_749_  (.B(\i_ibex/id_stage_i/controller_i/_241_ ),
    .C(\i_ibex/id_stage_i/controller_i/_228_ ),
    .A(\i_ibex/id_stage_i/controller_i/_031_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_306_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/controller_i/_750_  (.A(\i_ibex/id_stage_i/controller_i/_249_ ),
    .B(\i_ibex/id_stage_i/controller_i/_255_ ),
    .C(\i_ibex/id_stage_i/controller_i/_287_ ),
    .D(\i_ibex/id_stage_i/controller_i/_306_ ),
    .X(\i_ibex/id_stage_i/controller_i/_307_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_751_  (.Y(\i_ibex/id_stage_i/controller_i/_308_ ),
    .A(\i_ibex/id_stage_i/controller_i/_276_ ),
    .B(\i_ibex/id_stage_i/controller_i/_307_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_752_  (.B1(\i_ibex/id_stage_i/controller_i/_308_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_309_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_298_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_305_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_753_  (.Y(\i_ibex/id_stage_i/controller_i/_001_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_303_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_309_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_298_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_276_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_754_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_310_ ),
    .A(net1486),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_755_  (.Y(\i_ibex/id_stage_i/controller_i/_311_ ),
    .B(\i_ibex/id_stage_i/controller_i/_044_ ),
    .A_N(\i_ibex/id_stage_i/controller_i/_213_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_756_  (.Y(\i_ibex/id_stage_i/controller_i/_312_ ),
    .A(\i_ibex/id_stage_i/controller_i/_260_ ),
    .B(\i_ibex/id_stage_i/controller_i/_311_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_757_  (.A(net1488),
    .B(\i_ibex/id_stage_i/controller_i/_263_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_758_  (.A(\i_ibex/id_stage_i/controller_i/_273_ ),
    .B(\i_ibex/id_stage_i/controller_i/_313_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_314_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/controller_i/_759_  (.A2(\i_ibex/id_stage_i/controller_i/_314_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_312_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_280_ ),
    .X(\i_ibex/id_stage_i/controller_i/_315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_760_  (.Y(\i_ibex/id_stage_i/controller_i/_316_ ),
    .A(\i_ibex/id_stage_i/controller_i/_310_ ),
    .B(\i_ibex/id_stage_i/controller_i/_307_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_761_  (.B1(\i_ibex/id_stage_i/controller_i/_316_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_317_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_298_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_305_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_762_  (.Y(\i_ibex/id_stage_i/controller_i/_002_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_315_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_317_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_298_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_763_  (.Y(\i_ibex/id_stage_i/controller_i/_318_ ),
    .A(\i_ibex/id_stage_i/controller_i/_258_ ),
    .B(\i_ibex/id_stage_i/controller_i/_311_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_764_  (.B1(\i_ibex/id_stage_i/controller_i/_268_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_319_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_242_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_256_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_765_  (.Y(\i_ibex/id_stage_i/controller_i/_320_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_319_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_272_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_318_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_766_  (.A(\i_ibex/id_stage_i/controller_i/_280_ ),
    .B(\i_ibex/id_stage_i/controller_i/_298_ ),
    .C(\i_ibex/id_stage_i/controller_i/_320_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_767_  (.A(net1486),
    .B(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ),
    .Y(\i_ibex/id_stage_i/controller_i/_321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_768_  (.Y(\i_ibex/id_stage_i/controller_i/_322_ ),
    .A(\i_ibex/id_stage_i/controller_i/_321_ ),
    .B(\i_ibex/id_stage_i/controller_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_769_  (.A(\i_ibex/id_stage_i/controller_i/_239_ ),
    .B(\i_ibex/id_stage_i/controller_i/_322_ ),
    .Y(\i_ibex/debug_cause [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/controller_i/_770_  (.A(\i_ibex/id_stage_i/controller_i/_322_ ),
    .B_N(\i_ibex/id_stage_i/controller_i/_239_ ),
    .Y(\i_ibex/debug_cause [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_771_  (.Y(\i_ibex/id_stage_i/controller_i/_323_ ),
    .B(net1738),
    .A_N(\i_ibex/trigger_match ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_772_  (.B(\i_ibex/id_stage_i/controller_i/_266_ ),
    .C(\i_ibex/id_stage_i/controller_i/_323_ ),
    .A(\i_ibex/id_stage_i/controller_i/_321_ ),
    .Y(\i_ibex/debug_cause [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_773_  (.B1(net1489),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_324_ ),
    .VSS(VSS),
    .A1(net1487),
    .A2(\i_ibex/id_stage_i/controller_i/_225_ ));
 sg13g2_and2_2 \i_ibex/id_stage_i/controller_i/_774_  (.A(\i_ibex/id_stage_i/controller_i/_215_ ),
    .B(\i_ibex/id_stage_i/controller_i/_324_ ),
    .X(\i_ibex/debug_csr_save ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_775_  (.B(\i_ibex/id_stage_i/controller_i/_218_ ),
    .C(\i_ibex/id_stage_i/controller_i/_215_ ),
    .A(net1448),
    .Y(\i_ibex/id_stage_i/controller_i/_325_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_776_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_207_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_325_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_004_ ),
    .B1(\i_ibex/csr_restore_dret_id ));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_777_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_326_ ),
    .A(\i_ibex/id_stage_i/controller_i/do_single_step_q ),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_778_  (.B(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .C(\i_ibex/debug_single_step ),
    .A(net704),
    .Y(\i_ibex/id_stage_i/controller_i/_327_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_779_  (.B1(\i_ibex/id_stage_i/controller_i/_327_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/do_single_step_d ),
    .VSS(VSS),
    .A1(net706),
    .A2(\i_ibex/id_stage_i/controller_i/_326_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_780_  (.B1(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_328_ ),
    .VSS(VSS),
    .A1(net1738),
    .A2(\i_ibex/id_stage_i/controller_i/_269_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_781_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_d ),
    .A(\i_ibex/id_stage_i/controller_i/_328_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_782_  (.VDD(VDD),
    .Y(\i_ibex/exc_cause [6]),
    .A(\i_ibex/id_stage_i/controller_i/_229_ ),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/controller_i/_783_  (.X(\i_ibex/exc_cause [5]),
    .A(\i_ibex/id_stage_i/controller_i/handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .B(net39),
    .C(\i_ibex/exc_cause [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_784_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_329_ ),
    .B(\i_ibex/irqs [9]),
    .A(\i_ibex/irqs [8]));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_785_  (.A(\i_ibex/irqs [10]),
    .B(\i_ibex/irqs [11]),
    .C(\i_ibex/id_stage_i/controller_i/_329_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/id_stage_i/controller_i/_786_  (.A(\i_ibex/irqs [14]),
    .B(\i_ibex/irqs [15]),
    .C(\i_ibex/irqs [12]),
    .Y(\i_ibex/id_stage_i/controller_i/_331_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/irqs [13]));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_787_  (.A(\i_ibex/irqs [6]),
    .B(\i_ibex/irqs [7]),
    .Y(\i_ibex/id_stage_i/controller_i/_332_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_788_  (.A(\i_ibex/irqs [4]),
    .B(\i_ibex/irqs [5]),
    .Y(\i_ibex/id_stage_i/controller_i/_333_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_789_  (.A(\i_ibex/id_stage_i/controller_i/_332_ ),
    .B(\i_ibex/id_stage_i/controller_i/_333_ ),
    .X(\i_ibex/id_stage_i/controller_i/_334_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_790_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_335_ ),
    .B(\i_ibex/irqs [3]),
    .A(\i_ibex/irqs [2]));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_791_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_336_ ),
    .B(\i_ibex/irqs [1]),
    .A(\i_ibex/irqs [0]));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_792_  (.A(\i_ibex/id_stage_i/controller_i/_335_ ),
    .B(\i_ibex/id_stage_i/controller_i/_336_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_337_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_793_  (.B(\i_ibex/id_stage_i/controller_i/_331_ ),
    .C(\i_ibex/id_stage_i/controller_i/_334_ ),
    .A(\i_ibex/id_stage_i/controller_i/_330_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_338_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_337_ ));
 sg13g2_a21oi_2 \i_ibex/id_stage_i/controller_i/_794_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/id_stage_i/controller_i/_229_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_339_ ),
    .A2(net40),
    .A1(\i_ibex/id_stage_i/controller_i/handle_irq_$_AND__Y_A_$_AND__Y_B ));
 sg13g2_and2_2 \i_ibex/id_stage_i/controller_i/_795_  (.A(\i_ibex/id_stage_i/controller_i/_338_ ),
    .B(\i_ibex/id_stage_i/controller_i/_339_ ),
    .X(\i_ibex/exc_cause [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_796_  (.Y(\i_ibex/id_stage_i/controller_i/_340_ ),
    .A(\i_ibex/id_stage_i/controller_i/_337_ ),
    .B(\i_ibex/id_stage_i/controller_i/_339_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_797_  (.Y(\i_ibex/id_stage_i/controller_i/_341_ ),
    .B(\i_ibex/id_stage_i/controller_i/_331_ ),
    .A_N(\i_ibex/irqs [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/controller_i/_798_  (.A(\i_ibex/irqs [10]),
    .B(\i_ibex/irqs [11]),
    .C(\i_ibex/id_stage_i/controller_i/_329_ ),
    .D(\i_ibex/id_stage_i/controller_i/_341_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_342_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_799_  (.Y(\i_ibex/id_stage_i/controller_i/_343_ ),
    .B(\i_ibex/id_stage_i/controller_i/_334_ ),
    .A_N(\i_ibex/id_stage_i/controller_i/_342_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_800_  (.B(\i_ibex/id_stage_i/controller_i/_119_ ),
    .C(\i_ibex/id_stage_i/controller_i/_205_ ),
    .A(\i_ibex/id_stage_i/ecall_insn_dec ),
    .Y(\i_ibex/id_stage_i/controller_i/_344_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_801_  (.B1(\i_ibex/id_stage_i/controller_i/_344_ ),
    .VDD(VDD),
    .Y(\i_ibex/exc_cause [3]),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_340_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_343_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_802_  (.B1(\i_ibex/id_stage_i/controller_i/_331_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_345_ ),
    .VSS(VSS),
    .A1(\i_ibex/irqs [16]),
    .A2(\i_ibex/irqs [18]));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_803_  (.Y(\i_ibex/id_stage_i/controller_i/_346_ ),
    .A(\i_ibex/id_stage_i/controller_i/_330_ ),
    .B(\i_ibex/id_stage_i/controller_i/_345_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_804_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_334_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_346_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_347_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_340_ ));
 sg13g2_a21o_2 \i_ibex/id_stage_i/controller_i/_805_  (.A2(net612),
    .A1(\i_ibex/id_stage_i/controller_i/_119_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_347_ ),
    .X(\i_ibex/exc_cause [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_806_  (.A(\i_ibex/irqs [14]),
    .B(\i_ibex/irqs [15]),
    .Y(\i_ibex/id_stage_i/controller_i/_348_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_807_  (.A(\i_ibex/irqs [12]),
    .B(\i_ibex/irqs [13]),
    .C(\i_ibex/id_stage_i/controller_i/_348_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_349_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_808_  (.A(\i_ibex/irqs [10]),
    .B(\i_ibex/irqs [11]),
    .C(\i_ibex/id_stage_i/controller_i/_349_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_350_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_809_  (.B1(\i_ibex/id_stage_i/controller_i/_332_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_351_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_329_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_350_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_810_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_333_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_351_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_352_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_335_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_811_  (.B1(\i_ibex/id_stage_i/controller_i/_338_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_353_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_336_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_352_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_812_  (.A(\i_ibex/id_stage_i/controller_i/illegal_insn_q ),
    .B(\i_ibex/id_stage_i/controller_i/_033_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_354_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_813_  (.B(\i_ibex/id_stage_i/ebrk_insn ),
    .C(\i_ibex/id_stage_i/controller_i/_224_ ),
    .A(\i_ibex/id_stage_i/controller_i/_207_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_355_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_814_  (.Y(\i_ibex/id_stage_i/controller_i/_356_ ),
    .A(\i_ibex/id_stage_i/ecall_insn_dec ),
    .B(\i_ibex/id_stage_i/controller_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_815_  (.B1(\i_ibex/id_stage_i/controller_i/_356_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_357_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/ecall_insn_dec ),
    .A2(\i_ibex/id_stage_i/controller_i/_355_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_816_  (.A(\i_ibex/id_stage_i/controller_i/_205_ ),
    .B(\i_ibex/id_stage_i/controller_i/_357_ ),
    .X(\i_ibex/id_stage_i/controller_i/_358_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_817_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_359_ ),
    .A(\i_ibex/id_stage_i/controller_i/_358_ ),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_818_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_360_ ),
    .B(\i_ibex/id_stage_i/ecall_insn_dec ),
    .A(\i_ibex/id_stage_i/ebrk_insn ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_819_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_036_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_360_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_361_ ),
    .B1(\i_ibex/instr_fetch_err ));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_820_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_362_ ),
    .B(\i_ibex/id_stage_i/controller_i/store_err_q ),
    .A(\i_ibex/id_stage_i/controller_i/illegal_insn_q ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_821_  (.B1(\i_ibex/id_stage_i/controller_i/_362_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_363_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_031_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_361_ ));
 sg13g2_a221oi_1 \i_ibex/id_stage_i/controller_i/_822_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/id_stage_i/controller_i/_363_ ),
    .C1(net1406),
    .B1(\i_ibex/id_stage_i/controller_i/_359_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_030_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_364_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_354_ ));
 sg13g2_a21o_2 \i_ibex/id_stage_i/controller_i/_823_  (.A2(\i_ibex/id_stage_i/controller_i/_353_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_339_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_364_ ),
    .X(\i_ibex/exc_cause [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/controller_i/_824_  (.A(\i_ibex/id_stage_i/controller_i/_354_ ),
    .B(net1454),
    .C(\i_ibex/id_stage_i/controller_i/_358_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_365_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_825_  (.B1(\i_ibex/id_stage_i/controller_i/exc_req_q ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_366_ ),
    .VSS(VSS),
    .A1(net1485),
    .A2(\i_ibex/id_stage_i/controller_i/_033_ ));
 sg13g2_a21o_1 \i_ibex/id_stage_i/controller_i/_826_  (.A2(\i_ibex/id_stage_i/controller_i/_366_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_030_ ),
    .B1(net1449),
    .X(\i_ibex/id_stage_i/controller_i/_367_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_827_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_368_ ),
    .A(\i_ibex/irqs [5]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_828_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/irqs [6]),
    .A2(\i_ibex/id_stage_i/controller_i/_368_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_369_ ),
    .B1(\i_ibex/irqs [4]));
 sg13g2_nor2_1 \i_ibex/id_stage_i/controller_i/_829_  (.A(\i_ibex/irqs [3]),
    .B(\i_ibex/id_stage_i/controller_i/_369_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_370_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_830_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_371_ ),
    .A(\i_ibex/irqs [9]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_831_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_372_ ),
    .A(\i_ibex/irqs [13]),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_832_  (.Y(\i_ibex/id_stage_i/controller_i/_373_ ),
    .B(\i_ibex/irqs [15]),
    .A_N(\i_ibex/irqs [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_833_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_372_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_373_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_374_ ),
    .B1(\i_ibex/irqs [12]));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_834_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_375_ ),
    .A(\i_ibex/irqs [10]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_835_  (.B1(\i_ibex/id_stage_i/controller_i/_375_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_376_ ),
    .VSS(VSS),
    .A1(\i_ibex/irqs [11]),
    .A2(\i_ibex/id_stage_i/controller_i/_374_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_836_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/controller_i/_371_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_376_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_377_ ),
    .B1(\i_ibex/irqs [8]));
 sg13g2_nor4_1 \i_ibex/id_stage_i/controller_i/_837_  (.A(\i_ibex/irqs [7]),
    .B(\i_ibex/irqs [5]),
    .C(\i_ibex/irqs [3]),
    .D(\i_ibex/id_stage_i/controller_i/_377_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_378_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/controller_i/_838_  (.A(\i_ibex/irqs [2]),
    .B(\i_ibex/irqs [0]),
    .C(\i_ibex/id_stage_i/controller_i/_370_ ),
    .D(\i_ibex/id_stage_i/controller_i/_378_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_379_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_839_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_380_ ),
    .A(\i_ibex/irqs [1]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_840_  (.B1(\i_ibex/id_stage_i/controller_i/_338_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_381_ ),
    .VSS(VSS),
    .A1(\i_ibex/irqs [0]),
    .A2(\i_ibex/id_stage_i/controller_i/_380_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_841_  (.B1(\i_ibex/id_stage_i/controller_i/_339_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_382_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_379_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_381_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_842_  (.B1(\i_ibex/id_stage_i/controller_i/_382_ ),
    .VDD(VDD),
    .Y(\i_ibex/exc_cause [0]),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_365_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_367_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_843_  (.Y(\i_ibex/id_stage_i/controller_i/_383_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_218_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_215_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_119_ ),
    .A1(\i_ibex/debug_mode ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_844_  (.VDD(VDD),
    .Y(\i_ibex/exc_pc_mux_id [1]),
    .A(\i_ibex/id_stage_i/controller_i/_383_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_845_  (.B1(\i_ibex/id_stage_i/controller_i/_325_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_384_ ),
    .VSS(VSS),
    .A1(\i_ibex/debug_mode ),
    .A2(net1406));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_846_  (.VDD(VDD),
    .Y(\i_ibex/exc_pc_mux_id [0]),
    .A(\i_ibex/id_stage_i/controller_i/_384_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_847_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/exc_req_d ),
    .A(\i_ibex/id_stage_i/controller_i/_255_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_848_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_385_ ),
    .A(\i_ibex/id_stage_i/controller_i/_311_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_849_  (.B1(\i_ibex/id_stage_i/controller_i/_218_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_386_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_215_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_238_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_850_  (.B1(\i_ibex/id_stage_i/controller_i/_386_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/flush_id ),
    .VSS(VSS),
    .A1(net1448),
    .A2(\i_ibex/id_stage_i/controller_i/_385_ ));
 sg13g2_a21o_1 \i_ibex/id_stage_i/controller_i/_851_  (.A2(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ),
    .A1(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .B1(net1487),
    .X(\i_ibex/id_stage_i/controller_i/_387_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_852_  (.B1(\i_ibex/id_stage_i/controller_i/_387_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_388_ ),
    .VSS(VSS),
    .A1(net1489),
    .A2(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_853_  (.B(\i_ibex/id_stage_i/controller_i/_310_ ),
    .C(\i_ibex/id_stage_i/controller_i/_388_ ),
    .A(\i_ibex/id_stage_i/controller_i/_276_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_389_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/controller_i/_854_  (.B(\i_ibex/id_stage_i/controller_i/_218_ ),
    .C(\i_ibex/id_stage_i/controller_i/_262_ ),
    .A(\i_ibex/id_stage_i/controller_i/_265_ ),
    .Y(\i_ibex/id_stage_i/controller_i/_390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/controller_i/_855_  (.Y(\i_ibex/instr_req_gated ),
    .A(\i_ibex/id_stage_i/controller_i/_389_ ),
    .B(\i_ibex/id_stage_i/controller_i/_390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/controller_i/_856_  (.A2(\i_ibex/id_stage_i/controller_i/_289_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_285_ ),
    .B1(\i_ibex/id_stage_i/flush_id ),
    .X(\i_ibex/instr_valid_clear ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/controller_i/_857_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_391_ ),
    .A(\i_ibex/nmi_mode ),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_858_  (.B(\i_ibex/id_stage_i/controller_i/handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .C(net41),
    .A(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .Y(\i_ibex/id_stage_i/controller_i/_392_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net1448));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_859_  (.B1(\i_ibex/id_stage_i/controller_i/_392_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_393_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_391_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_228_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_860_  (.Y(\i_ibex/id_stage_i/controller_i/_394_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_217_ ),
    .B2(\i_ibex/id_stage_i/controller_i/_393_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_204_ ),
    .A1(\i_ibex/nmi_mode ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_861_  (.B1(\i_ibex/id_stage_i/controller_i/_394_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_005_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_391_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_042_ ));
 sg13g2_nor4_2 \i_ibex/id_stage_i/controller_i/_862_  (.A(\i_ibex/id_stage_i/controller_i/_201_ ),
    .B(\i_ibex/id_stage_i/mret_insn_dec ),
    .C(net1448),
    .Y(\i_ibex/pc_mux_id [2]),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_202_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/controller_i/_863_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net704),
    .A2(\i_ibex/id_stage_i/mret_insn_dec ),
    .Y(\i_ibex/id_stage_i/controller_i/_395_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_044_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_864_  (.B1(\i_ibex/id_stage_i/controller_i/_219_ ),
    .VDD(VDD),
    .Y(\i_ibex/pc_mux_id [1]),
    .VSS(VSS),
    .A1(net1448),
    .A2(\i_ibex/id_stage_i/controller_i/_395_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/controller_i/_865_  (.Y(\i_ibex/pc_mux_id [0]),
    .B(\i_ibex/id_stage_i/controller_i/_204_ ),
    .A_N(net694),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_866_  (.Y(\i_ibex/id_stage_i/controller_i/_396_ ),
    .A(\i_ibex/id_stage_i/controller_i/_044_ ),
    .B(\i_ibex/id_stage_i/controller_i/_213_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/controller_i/_867_  (.B1(\i_ibex/id_stage_i/controller_i/_396_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/controller_i/_397_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/controller_i/_202_ ),
    .A2(\i_ibex/id_stage_i/controller_i/_247_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/controller_i/_868_  (.Y(\i_ibex/id_stage_i/controller_i/_398_ ),
    .A(\i_ibex/id_stage_i/controller_i/_042_ ),
    .B(\i_ibex/id_stage_i/controller_i/_397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/controller_i/_869_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/controller_i/_399_ ),
    .B(\i_ibex/id_stage_i/jump_set ),
    .A(\i_ibex/id_stage_i/branch_set ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/controller_i/_870_  (.Y(\i_ibex/id_stage_i/controller_i/_400_ ),
    .B1(\i_ibex/id_stage_i/controller_i/_399_ ),
    .B2(net694),
    .A2(\i_ibex/id_stage_i/controller_i/_266_ ),
    .A1(\i_ibex/id_stage_i/controller_i/_261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/controller_i/_871_  (.B(\i_ibex/id_stage_i/controller_i/_389_ ),
    .C(\i_ibex/id_stage_i/controller_i/_398_ ),
    .A(\i_ibex/id_stage_i/controller_i/_229_ ),
    .Y(\i_ibex/pc_set ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/controller_i/_400_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_872_  (.A(\i_ibex/id_stage_i/jump_set ),
    .B(\i_ibex/id_stage_i/controller_run ),
    .X(\i_ibex/perf_jump ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/controller_i/_873_  (.A(\i_ibex/id_stage_i/branch_set ),
    .B(\i_ibex/id_stage_i/controller_run ),
    .X(\i_ibex/perf_tbranch ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/ctrl_fsm_cs[0]_reg  (.CLK(clknet_leaf_87_clk_i_regs),
    .RESET_B(net1611),
    .D(\i_ibex/id_stage_i/controller_i/_000_ ),
    .Q_N(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A ),
    .Q(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/id_stage_i/controller_i/ctrl_fsm_cs[1]_reg  (.RESET_B(net1611),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/id_stage_i/controller_i/_001_ ),
    .Q(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [1]),
    .Q_N(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_86_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/ctrl_fsm_cs[2]_reg  (.CLK(clknet_leaf_85_clk_i_regs),
    .RESET_B(net1610),
    .D(\i_ibex/id_stage_i/controller_i/_002_ ),
    .Q_N(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__B_Y_$_OR__Y_A ),
    .Q(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/id_stage_i/controller_i/ctrl_fsm_cs[3]_reg  (.RESET_B(net1610),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/id_stage_i/controller_i/_003_ ),
    .Q(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [3]),
    .Q_N(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__Y_B ),
    .CLK(clknet_leaf_85_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/id_stage_i/controller_i/debug_mode_o_reg  (.RESET_B(net1611),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/id_stage_i/controller_i/_004_ ),
    .Q(\i_ibex/debug_mode ),
    .Q_N(\i_ibex/id_stage_i/controller_i/debug_mode_o_$_NOT__A_Y ),
    .CLK(clknet_leaf_84_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/do_single_step_q_reg  (.CLK(clknet_leaf_85_clk_i_regs),
    .RESET_B(net1611),
    .D(\i_ibex/id_stage_i/controller_i/do_single_step_d ),
    .Q_N(\i_ibex/id_stage_i/controller_i/_403_ ),
    .Q(\i_ibex/id_stage_i/controller_i/do_single_step_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_q_reg  (.CLK(clknet_leaf_86_clk_i_regs),
    .RESET_B(net1610),
    .D(\i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_d ),
    .Q_N(\i_ibex/id_stage_i/controller_i/_404_ ),
    .Q(\i_ibex/id_stage_i/controller_i/enter_debug_mode_prio_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/exc_req_q_reg  (.CLK(clknet_leaf_87_clk_i_regs),
    .RESET_B(net1577),
    .D(\i_ibex/id_stage_i/controller_i/exc_req_d ),
    .Q_N(\i_ibex/id_stage_i/controller_i/_405_ ),
    .Q(\i_ibex/id_stage_i/controller_i/exc_req_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/illegal_insn_q_reg  (.CLK(clknet_leaf_88_clk_i_regs),
    .RESET_B(net1576),
    .D(\i_ibex/id_stage_i/controller_i/illegal_insn_d ),
    .Q_N(\i_ibex/id_stage_i/controller_i/_406_ ),
    .Q(\i_ibex/id_stage_i/controller_i/illegal_insn_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/load_err_q_reg  (.CLK(clknet_leaf_89_clk_i_regs),
    .RESET_B(net1577),
    .D(\i_ibex/lsu_load_err ),
    .Q_N(\i_ibex/id_stage_i/controller_i/_402_ ),
    .Q(\i_ibex/id_stage_i/controller_i/load_err_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/id_stage_i/controller_i/nmi_mode_o_reg  (.RESET_B(net1611),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/id_stage_i/controller_i/_005_ ),
    .Q(\i_ibex/nmi_mode ),
    .Q_N(\i_ibex/id_stage_i/controller_i/handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .CLK(clknet_leaf_84_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/controller_i/store_err_q_reg  (.CLK(clknet_leaf_89_clk_i_regs),
    .RESET_B(net1576),
    .D(\i_ibex/lsu_store_err ),
    .Q_N(\i_ibex/id_stage_i/controller_i/_401_ ),
    .Q(\i_ibex/id_stage_i/controller_i/store_err_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/decoder_i/_238_  (.Y(\i_ibex/id_stage_i/decoder_i/_227_ ),
    .A(\i_ibex/instr_rdata_id [0]),
    .B(\i_ibex/instr_rdata_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout600 (.A(net605),
    .X(net600),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_244_  (.A(\i_ibex/instr_rdata_id [0]),
    .B(\i_ibex/instr_rdata_id [1]),
    .X(\i_ibex/id_stage_i/decoder_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_245_  (.A(net719),
    .B(net738),
    .Y(\i_ibex/id_stage_i/decoder_i/_234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/id_stage_i/decoder_i/_246_  (.X(\i_ibex/id_stage_i/decoder_i/_235_ ),
    .A(net712),
    .B(\i_ibex/id_stage_i/decoder_i/_233_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_234_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/decoder_i/_247_  (.A(net772),
    .B(net709),
    .C(net715),
    .D(\i_ibex/id_stage_i/decoder_i/_235_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_236_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_249_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_001_ ),
    .A(net708),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_250_  (.A(\i_ibex/id_stage_i/decoder_i/_001_ ),
    .B(net715),
    .Y(\i_ibex/id_stage_i/decoder_i/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/decoder_i/_251_  (.A2(\i_ibex/id_stage_i/decoder_i/_002_ ),
    .A1(net740),
    .B1(\i_ibex/id_stage_i/decoder_i/_234_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout594 (.A(\i_ibex/alu_operand_a_ex [23]),
    .X(net594),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_253_  (.A(net717),
    .B_N(net739),
    .Y(\i_ibex/id_stage_i/decoder_i/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_254_  (.A(net721),
    .B_N(net715),
    .Y(\i_ibex/id_stage_i/decoder_i/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_255_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net721),
    .A2(\i_ibex/id_stage_i/decoder_i/_005_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_007_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_006_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_256_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_008_ ),
    .B(net739),
    .A(net721));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_257_  (.B1(\i_ibex/id_stage_i/decoder_i/_008_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_009_ ),
    .VSS(VSS),
    .A1(net713),
    .A2(\i_ibex/id_stage_i/decoder_i/_007_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_258_  (.Y(\i_ibex/id_stage_i/decoder_i/_010_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_009_ ),
    .B2(\i_ibex/id_stage_i/decoder_i/_001_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_003_ ),
    .A1(net712),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_259_  (.A(\i_ibex/id_stage_i/decoder_i/_227_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_236_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_010_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_260_  (.B(net739),
    .C(\i_ibex/instr_rdata_id [0]),
    .A(net720),
    .Y(\i_ibex/id_stage_i/decoder_i/_012_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/instr_rdata_id [1]));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_261_  (.A(net717),
    .B(\i_ibex/id_stage_i/decoder_i/_012_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout592 (.A(\i_ibex/alu_operand_a_ex [22]),
    .X(net592),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_264_  (.A(net772),
    .B(net780),
    .C(net776),
    .Y(\i_ibex/id_stage_i/decoder_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_265_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_017_ ),
    .B(net713),
    .A(net708));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_266_  (.Y(\i_ibex/id_stage_i/decoder_i/_018_ ),
    .A(net711),
    .B(net712),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_267_  (.B1(\i_ibex/id_stage_i/decoder_i/_018_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_019_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_016_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_017_ ));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_269_  (.A(net697),
    .B_N(net713),
    .Y(\i_ibex/id_stage_i/decoder_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_270_  (.A(net708),
    .B(net712),
    .Y(\i_ibex/id_stage_i/decoder_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_271_  (.A(net738),
    .B(\i_ibex/id_stage_i/decoder_i/_022_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_272_  (.Y(\i_ibex/id_stage_i/decoder_i/_024_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_023_ ),
    .B2(net718),
    .A2(\i_ibex/id_stage_i/decoder_i/_021_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_273_  (.A(net720),
    .B(\i_ibex/id_stage_i/decoder_i/_227_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_024_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_274_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_013_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_019_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_026_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_025_ ));
 sg13g2_nand2_2 \i_ibex/id_stage_i/decoder_i/_275_  (.Y(\i_ibex/id_stage_i/alu_op_a_mux_sel_dec [1]),
    .A(\i_ibex/id_stage_i/decoder_i/_011_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_276_  (.A(net771),
    .B(net776),
    .Y(\i_ibex/id_stage_i/decoder_i/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_277_  (.A(net717),
    .B(\i_ibex/id_stage_i/decoder_i/_012_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_027_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_017_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/id_stage_i/decoder_i/_278_  (.Y(\i_ibex/id_stage_i/alu_op_a_mux_sel_dec [0]),
    .B(\i_ibex/id_stage_i/decoder_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/decoder_i/_028_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_279_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_029_ ),
    .B(net716),
    .A(net771));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_280_  (.Y(\i_ibex/id_stage_i/decoder_i/_030_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_029_ ),
    .B2(\i_ibex/id_stage_i/decoder_i/_001_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_002_ ),
    .A1(net697),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/id_stage_i/decoder_i/_281_  (.Y(\i_ibex/id_stage_i/alu_op_b_mux_sel_dec ),
    .B(\i_ibex/id_stage_i/decoder_i/_235_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/decoder_i/_030_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_282_  (.A(net738),
    .B(net708),
    .X(\i_ibex/id_stage_i/decoder_i/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_283_  (.B1(net712),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_032_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_234_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_031_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_284_  (.B(net739),
    .C(\i_ibex/id_stage_i/decoder_i/_022_ ),
    .A(net720),
    .Y(\i_ibex/id_stage_i/decoder_i/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_285_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_032_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_033_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_034_ ),
    .B1(net715));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_286_  (.A(net720),
    .B(net708),
    .C(\i_ibex/id_stage_i/decoder_i/_005_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_287_  (.B1(\i_ibex/id_stage_i/decoder_i/_233_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_036_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_034_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_035_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_288_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_037_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_036_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_028_ ));
 sg13g2_xor2_1 \i_ibex/id_stage_i/decoder_i/_289_  (.B(net780),
    .A(net771),
    .X(\i_ibex/id_stage_i/decoder_i/_038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout590 (.A(\i_ibex/csr_addr [2]),
    .X(net590),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_291_  (.B1(net736),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_040_ ),
    .VSS(VSS),
    .A1(net750),
    .A2(\i_ibex/id_stage_i/decoder_i/_038_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_292_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_041_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_040_ ),
    .VSS(VSS));
 sg13g2_or4_2 \i_ibex/id_stage_i/decoder_i/_293_  (.A(net731),
    .B(net741),
    .C(net745),
    .D(net743),
    .X(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_294_  (.A(net748),
    .B(\i_ibex/id_stage_i/decoder_i/_041_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_295_  (.A(net770),
    .B(net750),
    .Y(\i_ibex/id_stage_i/decoder_i/_044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_296_  (.B1(net776),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_045_ ),
    .VSS(VSS),
    .A1(net736),
    .A2(\i_ibex/id_stage_i/decoder_i/_044_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_297_  (.A(net710),
    .B_N(net716),
    .Y(\i_ibex/id_stage_i/decoder_i/_046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_298_  (.Y(\i_ibex/id_stage_i/decoder_i/_047_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_235_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_299_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_043_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_045_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_048_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_047_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_300_  (.A(net715),
    .B(\i_ibex/id_stage_i/decoder_i/_018_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_301_  (.Y(\i_ibex/id_stage_i/decoder_i/_050_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_049_ ),
    .B2(net696),
    .A2(\i_ibex/id_stage_i/decoder_i/_022_ ),
    .A1(net715),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_302_  (.A(\i_ibex/id_stage_i/decoder_i/_227_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_008_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/decoder_i/_303_  (.B(\i_ibex/id_stage_i/decoder_i/_051_ ),
    .C(net775),
    .Y(\i_ibex/id_stage_i/decoder_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/decoder_i/_050_ ));
 sg13g2_nor2b_2 \i_ibex/id_stage_i/decoder_i/_304_  (.A(net776),
    .B_N(net778),
    .Y(\i_ibex/id_stage_i/decoder_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_305_  (.Y(\i_ibex/id_stage_i/decoder_i/_054_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_001_ ),
    .B(net716),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/id_stage_i/decoder_i/_306_  (.A(net713),
    .B(\i_ibex/id_stage_i/decoder_i/_227_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_008_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_055_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_054_ ));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_307_  (.B(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_053_ ),
    .A(net773),
    .Y(\i_ibex/id_stage_i/decoder_i/_056_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_055_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_308_  (.B1(\i_ibex/id_stage_i/decoder_i/_056_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_057_ ),
    .VSS(VSS),
    .A1(net771),
    .A2(\i_ibex/id_stage_i/decoder_i/_052_ ));
 sg13g2_or3_2 \i_ibex/id_stage_i/decoder_i/_309_  (.A(\i_ibex/id_stage_i/decoder_i/_037_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_048_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_057_ ),
    .X(\i_ibex/alu_operator_ex [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_310_  (.B(net696),
    .C(\i_ibex/id_stage_i/decoder_i/_002_ ),
    .A(net714),
    .Y(\i_ibex/id_stage_i/decoder_i/_058_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_051_ ));
 sg13g2_nor2b_2 \i_ibex/id_stage_i/decoder_i/_311_  (.A(net773),
    .B_N(net774),
    .Y(\i_ibex/id_stage_i/decoder_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_312_  (.A(\i_ibex/id_stage_i/decoder_i/_058_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_059_ ),
    .Y(\i_ibex/alu_operator_ex [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_313_  (.A(net748),
    .B(\i_ibex/id_stage_i/decoder_i/_053_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_059_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_060_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_314_  (.B1(net736),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_061_ ),
    .VSS(VSS),
    .A1(net770),
    .A2(net751));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_315_  (.A(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .B_N(\i_ibex/id_stage_i/decoder_i/_061_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_316_  (.B1(\i_ibex/id_stage_i/decoder_i/_062_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_063_ ),
    .VSS(VSS),
    .A1(net751),
    .A2(\i_ibex/id_stage_i/decoder_i/_060_ ));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_317_  (.Y(\i_ibex/id_stage_i/decoder_i/_064_ ),
    .B(net736),
    .A_N(net770),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_318_  (.A(net736),
    .B(net780),
    .Y(\i_ibex/id_stage_i/decoder_i/_065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_319_  (.Y(\i_ibex/id_stage_i/decoder_i/_066_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_065_ ),
    .B2(\i_ibex/id_stage_i/decoder_i/_059_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_064_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_320_  (.A(net751),
    .B(net748),
    .C(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_067_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_321_  (.A(\i_ibex/id_stage_i/decoder_i/_066_ ),
    .B_N(\i_ibex/id_stage_i/decoder_i/_067_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_322_  (.A(net748),
    .B(\i_ibex/id_stage_i/decoder_i/_063_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_068_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_323_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_070_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_059_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_053_ ));
 sg13g2_and4_1 \i_ibex/id_stage_i/decoder_i/_324_  (.A(net713),
    .B(net696),
    .C(\i_ibex/id_stage_i/decoder_i/_002_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_051_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_325_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_055_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_070_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_072_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_071_ ));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_326_  (.B1(\i_ibex/id_stage_i/decoder_i/_072_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_073_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_047_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_069_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_327_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/alu_operator_ex [3]),
    .B(\i_ibex/id_stage_i/decoder_i/_073_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_037_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_328_  (.B(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_055_ ),
    .A(net773),
    .Y(\i_ibex/id_stage_i/decoder_i/_074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_329_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_075_ ),
    .A(net778),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_330_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_052_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_074_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_076_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_075_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_331_  (.A(net751),
    .B(\i_ibex/id_stage_i/decoder_i/_075_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_332_  (.B1(net776),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_078_ ),
    .VSS(VSS),
    .A1(net735),
    .A2(\i_ibex/id_stage_i/decoder_i/_077_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_333_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_043_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_078_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_079_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_047_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_334_  (.A(net771),
    .B(\i_ibex/id_stage_i/decoder_i/_058_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/id_stage_i/decoder_i/_335_  (.A(\i_ibex/id_stage_i/decoder_i/_037_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_076_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_079_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_080_ ),
    .X(\i_ibex/alu_operator_ex [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_336_  (.Y(\i_ibex/id_stage_i/decoder_i/_081_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_067_ ),
    .A_N(\i_ibex/id_stage_i/decoder_i/_066_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_337_  (.Y(\i_ibex/id_stage_i/decoder_i/_082_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_063_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_338_  (.A(\i_ibex/id_stage_i/decoder_i/_047_ ),
    .B_N(\i_ibex/id_stage_i/decoder_i/_067_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_083_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_339_  (.A(\i_ibex/id_stage_i/decoder_i/_075_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_027_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_340_  (.A(net735),
    .B(\i_ibex/id_stage_i/decoder_i/_016_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_084_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_085_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_341_  (.B(\i_ibex/id_stage_i/decoder_i/_083_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_085_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_082_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_342_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_087_ ),
    .A(net771),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_343_  (.Y(\i_ibex/id_stage_i/decoder_i/_088_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_075_ ),
    .B(net774),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_344_  (.Y(\i_ibex/id_stage_i/decoder_i/_089_ ),
    .B(net778),
    .A_N(net774),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_345_  (.B1(\i_ibex/id_stage_i/decoder_i/_089_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_090_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_087_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_088_ ));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_346_  (.Y(\i_ibex/id_stage_i/decoder_i/_091_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_087_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_347_  (.B1(\i_ibex/id_stage_i/decoder_i/_091_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_092_ ),
    .VSS(VSS),
    .A1(net778),
    .A2(\i_ibex/id_stage_i/decoder_i/_027_ ));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_348_  (.Y(\i_ibex/id_stage_i/decoder_i/_093_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_092_ ),
    .B2(\i_ibex/id_stage_i/decoder_i/_055_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_090_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_349_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_086_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_093_ ),
    .Y(\i_ibex/alu_operator_ex [1]),
    .B1(\i_ibex/id_stage_i/decoder_i/_036_ ));
 sg13g2_mux2_1 \i_ibex/id_stage_i/decoder_i/_350_  (.A0(\i_ibex/id_stage_i/decoder_i/_064_ ),
    .A1(net735),
    .S(net774),
    .X(\i_ibex/id_stage_i/decoder_i/_094_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/decoder_i/_351_  (.B(\i_ibex/id_stage_i/decoder_i/_053_ ),
    .C(net771),
    .Y(\i_ibex/id_stage_i/decoder_i/_095_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net735));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_352_  (.B1(\i_ibex/id_stage_i/decoder_i/_095_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_096_ ),
    .VSS(VSS),
    .A1(net778),
    .A2(\i_ibex/id_stage_i/decoder_i/_094_ ));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_353_  (.B(\i_ibex/id_stage_i/decoder_i/_083_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_096_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_043_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_354_  (.B1(\i_ibex/id_stage_i/decoder_i/_088_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_098_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_042_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_095_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_355_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_087_ ),
    .A2(net780),
    .Y(\i_ibex/id_stage_i/decoder_i/_099_ ),
    .B1(net774));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_356_  (.Y(\i_ibex/id_stage_i/decoder_i/_100_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_099_ ),
    .B2(\i_ibex/id_stage_i/decoder_i/_071_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_098_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_357_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_097_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_100_ ),
    .Y(\i_ibex/alu_operator_ex [0]),
    .B1(\i_ibex/id_stage_i/decoder_i/_036_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_358_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_101_ ),
    .B(net742),
    .A(net743));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_359_  (.A(net751),
    .B(net749),
    .C(net731),
    .D(net746),
    .Y(\i_ibex/id_stage_i/decoder_i/_102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_360_  (.A(\i_ibex/id_stage_i/decoder_i/_101_ ),
    .B_N(\i_ibex/id_stage_i/decoder_i/_102_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/id_stage_i/decoder_i/_362_  (.Y(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .A(net773),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_363_  (.Y(\i_ibex/id_stage_i/decoder_i/_106_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .B(net735),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout588 (.A(net590),
    .X(net588),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(net590),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(net590),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/id_stage_i/decoder_i/_367_  (.Y(\i_ibex/id_stage_i/decoder_i/_110_ ),
    .B(net779),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net775));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_368_  (.Y(\i_ibex/id_stage_i/decoder_i/_111_ ),
    .A(\i_ibex/instr_rdata_id [0]),
    .B(\i_ibex/instr_rdata_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_369_  (.A(net714),
    .B(net710),
    .C(\i_ibex/id_stage_i/decoder_i/_110_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_111_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_370_  (.A(net738),
    .B(net719),
    .Y(\i_ibex/id_stage_i/decoder_i/_113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_371_  (.B(\i_ibex/id_stage_i/decoder_i/_112_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_113_ ),
    .A(net717),
    .Y(\i_ibex/id_stage_i/decoder_i/_114_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_372_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_103_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_106_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_115_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_114_ ));
 sg13g2_buf_1 fanout585 (.A(\i_ibex/alu_operand_a_ex [31]),
    .X(net585),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_374_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_117_ ),
    .A(net710),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_375_  (.B1(net777),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_118_ ),
    .VSS(VSS),
    .A1(net708),
    .A2(net779));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_376_  (.A(net772),
    .B(\i_ibex/id_stage_i/decoder_i/_118_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_377_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_117_ ),
    .A2(\i_ibex/id_stage_i/imm_u_type [14]),
    .Y(\i_ibex/id_stage_i/decoder_i/_120_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_119_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_378_  (.A(\i_ibex/instr_rdata_id [0]),
    .B(\i_ibex/instr_rdata_id [1]),
    .X(\i_ibex/id_stage_i/decoder_i/_121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_379_  (.A(\i_ibex/id_stage_i/decoder_i/_121_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_113_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/id_stage_i/decoder_i/_380_  (.A(net717),
    .B_N(net714),
    .Y(\i_ibex/id_stage_i/decoder_i/_123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/decoder_i/_381_  (.Y(\i_ibex/id_stage_i/decoder_i/_124_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_122_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_382_  (.A(\i_ibex/id_stage_i/decoder_i/_120_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_124_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_383_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_126_ ),
    .A(net775),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_384_  (.Y(\i_ibex/id_stage_i/decoder_i/_127_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_126_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_385_  (.B(net719),
    .C(\i_ibex/id_stage_i/decoder_i/_127_ ),
    .A(net740),
    .Y(\i_ibex/id_stage_i/decoder_i/_128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_386_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_129_ ),
    .B(net779),
    .A(net772));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_387_  (.B(\i_ibex/id_stage_i/decoder_i/_113_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_129_ ),
    .A(net776),
    .Y(\i_ibex/id_stage_i/decoder_i/_130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/id_stage_i/decoder_i/_388_  (.A(net717),
    .B(net714),
    .C(net710),
    .D(\i_ibex/id_stage_i/decoder_i/_111_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_389_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_128_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_130_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_132_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_131_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_390_  (.A(net755),
    .B_N(net741),
    .Y(\i_ibex/id_stage_i/decoder_i/_133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_391_  (.A(net761),
    .B_N(net757),
    .Y(\i_ibex/id_stage_i/decoder_i/_134_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/decoder_i/_392_  (.A(net751),
    .B(net745),
    .C(net735),
    .D(net753),
    .X(\i_ibex/id_stage_i/decoder_i/_135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_393_  (.B(\i_ibex/id_stage_i/decoder_i/_133_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_134_ ),
    .A(net744),
    .Y(\i_ibex/id_stage_i/decoder_i/_136_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_135_ ));
 sg13g2_nor4_2 \i_ibex/id_stage_i/decoder_i/_394_  (.A(net751),
    .B(net746),
    .C(net735),
    .Y(\i_ibex/id_stage_i/decoder_i/_137_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/imm_u_type [24]));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_395_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_138_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_137_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_396_  (.B1(\i_ibex/id_stage_i/decoder_i/_138_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_139_ ),
    .VSS(VSS),
    .A1(net754),
    .A2(\i_ibex/id_stage_i/decoder_i/_136_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_397_  (.A(net768),
    .B(net766),
    .Y(\i_ibex/id_stage_i/decoder_i/_140_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_398_  (.A(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .B(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .C(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .Y(\i_ibex/id_stage_i/decoder_i/_141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_399_  (.Y(\i_ibex/id_stage_i/decoder_i/_142_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_140_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_400_  (.A(net748),
    .B(net731),
    .Y(\i_ibex/id_stage_i/decoder_i/_143_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_401_  (.A(net770),
    .B(net779),
    .C(\i_ibex/id_stage_i/imm_u_type [13]),
    .Y(\i_ibex/id_stage_i/decoder_i/_144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/decoder_i/_402_  (.B(\i_ibex/id_stage_i/decoder_i/_143_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_144_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_145_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net754));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_403_  (.A(\i_ibex/id_stage_i/imm_s_type [4]),
    .B(\i_ibex/id_stage_i/imm_s_type [3]),
    .Y(\i_ibex/id_stage_i/decoder_i/_146_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_404_  (.A(\i_ibex/id_stage_i/imm_s_type [2]),
    .B(\i_ibex/id_stage_i/imm_s_type [0]),
    .C(\i_ibex/id_stage_i/imm_s_type [1]),
    .Y(\i_ibex/id_stage_i/decoder_i/_147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_405_  (.Y(\i_ibex/id_stage_i/decoder_i/_148_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_146_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_406_  (.A(\i_ibex/id_stage_i/decoder_i/_142_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_145_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_148_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_149_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_407_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_150_ ),
    .B(net775),
    .A(net779));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_408_  (.A(net715),
    .B(net713),
    .X(\i_ibex/id_stage_i/decoder_i/_151_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_409_  (.B(\i_ibex/id_stage_i/decoder_i/_121_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_113_ ),
    .A(net710),
    .Y(\i_ibex/id_stage_i/decoder_i/_152_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_151_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_410_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_153_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_152_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_150_ ));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_411_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_139_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_149_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_154_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_153_ ));
 sg13g2_or4_2 \i_ibex/id_stage_i/decoder_i/_412_  (.A(\i_ibex/id_stage_i/decoder_i/_115_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_125_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_132_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_154_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout584 (.A(net585),
    .X(net584),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_414_  (.A(\i_ibex/id_stage_i/decoder_i/_133_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_134_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_415_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_158_ ),
    .A(net755),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_416_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_159_ ),
    .A(net761),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_417_  (.A(net741),
    .B(\i_ibex/id_stage_i/decoder_i/_158_ ),
    .C(net757),
    .D(\i_ibex/id_stage_i/decoder_i/_159_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_160_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_418_  (.B1(net744),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_161_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_157_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_160_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_419_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_162_ ),
    .A(net759),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/decoder_i/_420_  (.B(\i_ibex/id_stage_i/decoder_i/_162_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_158_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_163_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/decoder_i/_101_ ));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/decoder_i/_421_  (.B(\i_ibex/id_stage_i/decoder_i/_161_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_163_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_164_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/id_stage_i/decoder_i/_153_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_422_  (.A(net776),
    .B_N(net748),
    .Y(\i_ibex/id_stage_i/decoder_i/_165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_423_  (.B1(\i_ibex/id_stage_i/decoder_i/_150_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_166_ ),
    .VSS(VSS),
    .A1(net735),
    .A2(\i_ibex/id_stage_i/decoder_i/_165_ ));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_424_  (.A(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .B(net748),
    .C(\i_ibex/id_stage_i/decoder_i/_110_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/decoder_i/_425_  (.A2(\i_ibex/id_stage_i/decoder_i/_166_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_167_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/id_stage_i/decoder_i/_426_  (.A(net746),
    .B(net743),
    .C(net742),
    .Y(\i_ibex/id_stage_i/decoder_i/_169_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net737));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_427_  (.A(net752),
    .B_N(net772),
    .Y(\i_ibex/id_stage_i/decoder_i/_170_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_428_  (.B(\i_ibex/id_stage_i/decoder_i/_143_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_169_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_110_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_171_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_170_ ));
 sg13g2_and4_1 \i_ibex/id_stage_i/decoder_i/_429_  (.A(\i_ibex/id_stage_i/decoder_i/_117_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_121_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_113_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_151_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_172_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_430_  (.Y(\i_ibex/id_stage_i/decoder_i/_173_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_171_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_172_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/decoder_i/_431_  (.A2(\i_ibex/id_stage_i/decoder_i/_168_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_103_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_173_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_174_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_432_  (.Y(\i_ibex/id_stage_i/decoder_i/_175_ ),
    .B(net719),
    .A_N(net709),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_433_  (.Y(\i_ibex/id_stage_i/decoder_i/_176_ ),
    .A(net714),
    .B(net709),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_434_  (.B1(\i_ibex/id_stage_i/decoder_i/_176_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_177_ ),
    .VSS(VSS),
    .A1(net713),
    .A2(\i_ibex/id_stage_i/decoder_i/_175_ ));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_435_  (.A(net718),
    .B_N(net738),
    .Y(\i_ibex/id_stage_i/decoder_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_436_  (.A(net714),
    .B_N(net709),
    .Y(\i_ibex/id_stage_i/decoder_i/_179_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_437_  (.Y(\i_ibex/id_stage_i/decoder_i/_180_ ),
    .B(net716),
    .A_N(net709),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_438_  (.B1(\i_ibex/id_stage_i/decoder_i/_180_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_181_ ),
    .VSS(VSS),
    .A1(net739),
    .A2(\i_ibex/id_stage_i/decoder_i/_179_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_439_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_182_ ),
    .A(net719),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/id_stage_i/decoder_i/_440_  (.Y(\i_ibex/id_stage_i/decoder_i/_183_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_181_ ),
    .B2(\i_ibex/id_stage_i/decoder_i/_182_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_178_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_177_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_441_  (.B(net709),
    .C(\i_ibex/id_stage_i/decoder_i/_121_ ),
    .A(net740),
    .Y(\i_ibex/id_stage_i/decoder_i/_184_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_123_ ));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_442_  (.A(net719),
    .B(\i_ibex/id_stage_i/decoder_i/_144_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_184_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_443_  (.A(\i_ibex/illegal_c_insn_id ),
    .B(\i_ibex/id_stage_i/decoder_i/_111_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_183_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_185_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_186_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/id_stage_i/decoder_i/_444_  (.B(\i_ibex/id_stage_i/decoder_i/_174_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_186_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_164_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 \i_ibex/id_stage_i/decoder_i/_445_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/illegal_insn_dec ),
    .B(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_155_ ));
 sg13g2_nor4_2 \i_ibex/id_stage_i/decoder_i/_446_  (.A(\i_ibex/id_stage_i/decoder_i/_117_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_124_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .Y(\i_ibex/id_stage_i/branch_in_dec ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_187_ ));
 sg13g2_or2_1 \i_ibex/id_stage_i/decoder_i/_447_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/id_stage_i/decoder_i/_188_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_144_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_152_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_448_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/rf_wdata_sel ),
    .A(\i_ibex/id_stage_i/decoder_i/_188_ ),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_449_  (.A(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_188_ ),
    .Y(\i_ibex/csr_access ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_450_  (.Y(\i_ibex/id_stage_i/decoder_i/_189_ ),
    .A(net776),
    .B(\i_ibex/id_stage_i/decoder_i/_142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_451_  (.A(\i_ibex/id_stage_i/decoder_i/_152_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_189_ ),
    .Y(\i_ibex/csr_op [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_452_  (.B1(net780),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_190_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_126_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_142_ ));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_453_  (.A(\i_ibex/id_stage_i/decoder_i/_152_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_190_ ),
    .Y(\i_ibex/csr_op [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/id_stage_i/decoder_i/_454_  (.B(\i_ibex/id_stage_i/decoder_i/_117_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_122_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_191_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net716));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_455_  (.A(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_191_ ),
    .Y(\i_ibex/id_stage_i/lsu_req_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_456_  (.A(net713),
    .B(net773),
    .C(\i_ibex/id_stage_i/decoder_i/_191_ ),
    .Y(\i_ibex/lsu_sign_ext ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_457_  (.A(\i_ibex/id_stage_i/decoder_i/_150_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_191_ ),
    .Y(\i_ibex/lsu_type [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_458_  (.A(\i_ibex/id_stage_i/decoder_i/_110_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_191_ ),
    .Y(\i_ibex/lsu_type [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/id_stage_i/decoder_i/_459_  (.A(net709),
    .B(\i_ibex/id_stage_i/decoder_i/_124_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .Y(\i_ibex/lsu_we ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_187_ ));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_460_  (.A(\i_ibex/id_stage_i/decoder_i/_152_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_145_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_136_ ),
    .Y(\i_ibex/id_stage_i/dret_insn_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_461_  (.A(\i_ibex/id_stage_i/decoder_i/_152_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_145_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/id_stage_i/decoder_i/_462_  (.Y(\i_ibex/id_stage_i/decoder_i/_193_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_137_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_463_  (.A(\i_ibex/id_stage_i/decoder_i/_159_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_163_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_193_ ),
    .Y(\i_ibex/id_stage_i/ebrk_insn ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_464_  (.A(net763),
    .B(\i_ibex/id_stage_i/decoder_i/_163_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_193_ ),
    .Y(\i_ibex/id_stage_i/ecall_insn_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_465_  (.Y(\i_ibex/id_stage_i/decoder_i/_194_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_075_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_466_  (.B(net716),
    .C(\i_ibex/id_stage_i/decoder_i/_235_ ),
    .A(net710),
    .Y(\i_ibex/id_stage_i/imm_a_mux_sel ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_194_ ));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_467_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_195_ ),
    .A(net720),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/id_stage_i/decoder_i/_468_  (.X(\i_ibex/id_stage_i/decoder_i/_196_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_195_ ),
    .B(net739),
    .C(\i_ibex/id_stage_i/decoder_i/_046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_469_  (.B1(\i_ibex/id_stage_i/decoder_i/_233_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_197_ ),
    .VSS(VSS),
    .A1(\i_ibex/id_stage_i/decoder_i/_034_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_196_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_470_  (.A(net738),
    .B(\i_ibex/id_stage_i/decoder_i/_233_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_471_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_195_ ),
    .A2(net696),
    .Y(\i_ibex/id_stage_i/decoder_i/_199_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_018_ ));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_472_  (.A(net771),
    .B(\i_ibex/id_stage_i/decoder_i/_012_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_017_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_089_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_473_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_198_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_199_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_201_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_200_ ));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_474_  (.A(net716),
    .B(\i_ibex/id_stage_i/decoder_i/_197_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_201_ ),
    .Y(\i_ibex/id_stage_i/imm_b_mux_sel_dec [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_475_  (.A(net739),
    .B(net716),
    .C(net696),
    .D(\i_ibex/id_stage_i/decoder_i/_018_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_476_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net738),
    .A2(\i_ibex/id_stage_i/decoder_i/_046_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_203_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_202_ ));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_477_  (.A(net720),
    .B(\i_ibex/id_stage_i/decoder_i/_227_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_203_ ),
    .Y(\i_ibex/id_stage_i/imm_b_mux_sel_dec [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_478_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_204_ ),
    .A(net696),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_479_  (.A(net720),
    .B(\i_ibex/id_stage_i/decoder_i/_054_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/id_stage_i/decoder_i/_480_  (.A2(\i_ibex/id_stage_i/decoder_i/_049_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_204_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_205_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_206_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_481_  (.A(net712),
    .B(\i_ibex/id_stage_i/decoder_i/_012_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_089_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_482_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net712),
    .A2(\i_ibex/id_stage_i/decoder_i/_051_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_208_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_207_ ));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_483_  (.A(net708),
    .B(\i_ibex/id_stage_i/decoder_i/_029_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_208_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_484_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_198_ ),
    .A2(\i_ibex/id_stage_i/decoder_i/_206_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_210_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_209_ ));
 sg13g2_nor2_2 \i_ibex/id_stage_i/decoder_i/_485_  (.A(\i_ibex/id_stage_i/decoder_i/_197_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_210_ ),
    .Y(\i_ibex/id_stage_i/imm_b_mux_sel_dec [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_486_  (.B(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_112_ ),
    .A(net719),
    .Y(\i_ibex/id_stage_i/decoder_i/_211_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_178_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_487_  (.A(\i_ibex/id_stage_i/decoder_i/_184_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_211_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_212_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_488_  (.A(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_212_ ),
    .Y(\i_ibex/id_stage_i/jump_in_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/id_stage_i/decoder_i/_489_  (.A(\i_ibex/id_stage_i/decoder_i/_204_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_212_ ),
    .Y(\i_ibex/id_stage_i/jump_set_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 \i_ibex/id_stage_i/decoder_i/_490_  (.A(net743),
    .B(\i_ibex/id_stage_i/decoder_i/_137_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_157_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_192_ ),
    .X(\i_ibex/id_stage_i/mret_insn_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/id_stage_i/decoder_i/_491_  (.A(net751),
    .B(\i_ibex/id_stage_i/decoder_i/_143_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_169_ ),
    .D(\i_ibex/id_stage_i/decoder_i/_172_ ),
    .X(\i_ibex/id_stage_i/decoder_i/_213_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_492_  (.A(net770),
    .B(\i_ibex/id_stage_i/decoder_i/_213_ ),
    .X(\i_ibex/multdiv_operator_ex [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/id_stage_i/decoder_i/_493_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/id_stage_i/decoder_i/_105_ ),
    .A2(net780),
    .Y(\i_ibex/id_stage_i/decoder_i/_214_ ),
    .B1(net775));
 sg13g2_nor2b_1 \i_ibex/id_stage_i/decoder_i/_494_  (.A(\i_ibex/id_stage_i/decoder_i/_214_ ),
    .B_N(\i_ibex/id_stage_i/decoder_i/_213_ ),
    .Y(\i_ibex/multdiv_operator_ex [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_495_  (.Y(\i_ibex/id_stage_i/decoder_i/_215_ ),
    .B(net772),
    .A_N(net779),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_496_  (.B1(\i_ibex/id_stage_i/decoder_i/_215_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_216_ ),
    .VSS(VSS),
    .A1(net772),
    .A2(\i_ibex/id_stage_i/decoder_i/_110_ ));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_497_  (.A(\i_ibex/id_stage_i/decoder_i/_213_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_216_ ),
    .X(\i_ibex/multdiv_signed_mode_ex [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/id_stage_i/decoder_i/_498_  (.B(\i_ibex/id_stage_i/decoder_i/_127_ ),
    .A(net779),
    .X(\i_ibex/id_stage_i/decoder_i/_217_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/id_stage_i/decoder_i/_499_  (.A(\i_ibex/id_stage_i/decoder_i/_213_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_217_ ),
    .X(\i_ibex/multdiv_signed_mode_ex [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_500_  (.Y(\i_ibex/id_stage_i/decoder_i/_218_ ),
    .A(net711),
    .B(\i_ibex/id_stage_i/decoder_i/_123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_501_  (.B1(\i_ibex/id_stage_i/decoder_i/_218_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_219_ ),
    .VSS(VSS),
    .A1(net739),
    .A2(net709));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_502_  (.A(net720),
    .B(\i_ibex/id_stage_i/decoder_i/_111_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_220_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/id_stage_i/decoder_i/_503_  (.Y(\i_ibex/id_stage_i/decoder_i/_221_ ),
    .A(\i_ibex/id_stage_i/decoder_i/_219_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_220_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_504_  (.B1(\i_ibex/id_stage_i/decoder_i/_221_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/rf_ren_a_dec ),
    .VSS(VSS),
    .A1(net772),
    .A2(\i_ibex/id_stage_i/decoder_i/_188_ ));
 sg13g2_a21o_1 \i_ibex/id_stage_i/decoder_i/_505_  (.A2(\i_ibex/id_stage_i/decoder_i/_123_ ),
    .A1(\i_ibex/id_stage_i/decoder_i/_122_ ),
    .B1(\i_ibex/id_stage_i/decoder_i/_172_ ),
    .X(\i_ibex/id_stage_i/rf_ren_b_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/id_stage_i/decoder_i/_506_  (.Y(\i_ibex/id_stage_i/decoder_i/_222_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_220_ ),
    .A_N(\i_ibex/id_stage_i/decoder_i/_180_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/id_stage_i/decoder_i/_507_  (.B1(\i_ibex/id_stage_i/decoder_i/_222_ ),
    .VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_223_ ),
    .VSS(VSS),
    .A1(net696),
    .A2(\i_ibex/id_stage_i/decoder_i/_184_ ));
 sg13g2_nor2_1 \i_ibex/id_stage_i/decoder_i/_508_  (.A(net1365),
    .B(\i_ibex/id_stage_i/decoder_i/_223_ ),
    .Y(\i_ibex/id_stage_i/decoder_i/_224_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/id_stage_i/decoder_i/_509_  (.A(\i_ibex/id_stage_i/decoder_i/_155_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_187_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_224_ ),
    .Y(\i_ibex/id_stage_i/rf_we_dec ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/id_stage_i/decoder_i/_510_  (.VDD(VDD),
    .Y(\i_ibex/id_stage_i/decoder_i/_225_ ),
    .A(net742),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/id_stage_i/decoder_i/_511_  (.B(\i_ibex/id_stage_i/decoder_i/_225_ ),
    .C(net756),
    .A(net744),
    .Y(\i_ibex/id_stage_i/decoder_i/_226_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/id_stage_i/decoder_i/_162_ ));
 sg13g2_nor3_2 \i_ibex/id_stage_i/decoder_i/_512_  (.A(\i_ibex/id_stage_i/decoder_i/_159_ ),
    .B(\i_ibex/id_stage_i/decoder_i/_193_ ),
    .C(\i_ibex/id_stage_i/decoder_i/_226_ ),
    .Y(\i_ibex/perf_wfi_wait ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/if_stage_i/_798__380  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net380));
 sg13g2_dfrbp_2 \i_ibex/id_stage_i/id_fsm_q_reg  (.RESET_B(net1656),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/id_stage_i/_0000_ ),
    .Q(\i_ibex/id_stage_i/id_fsm_q ),
    .Q_N(\i_ibex/id_stage_i/instr_first_cycle_id_o_$_AND__Y_B ),
    .CLK(clknet_leaf_89_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[0]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1527),
    .D(\i_ibex/id_stage_i/_0001_ ),
    .Q_N(\i_ibex/id_stage_i/_0626_ ),
    .Q(\i_ibex/imd_val_q_ex [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[10]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0002_ ),
    .Q_N(\i_ibex/id_stage_i/_0625_ ),
    .Q(\i_ibex/imd_val_q_ex [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[11]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0003_ ),
    .Q_N(\i_ibex/id_stage_i/_0624_ ),
    .Q(\i_ibex/imd_val_q_ex [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[12]_reg  (.CLK(clknet_leaf_0_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0004_ ),
    .Q_N(\i_ibex/id_stage_i/_0623_ ),
    .Q(\i_ibex/imd_val_q_ex [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[13]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0005_ ),
    .Q_N(\i_ibex/id_stage_i/_0622_ ),
    .Q(\i_ibex/imd_val_q_ex [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[14]_reg  (.CLK(clknet_leaf_0_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0006_ ),
    .Q_N(\i_ibex/id_stage_i/_0621_ ),
    .Q(\i_ibex/imd_val_q_ex [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[15]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0007_ ),
    .Q_N(\i_ibex/id_stage_i/_0620_ ),
    .Q(\i_ibex/imd_val_q_ex [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[16]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0008_ ),
    .Q_N(\i_ibex/id_stage_i/_0619_ ),
    .Q(\i_ibex/imd_val_q_ex [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[17]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1527),
    .D(\i_ibex/id_stage_i/_0009_ ),
    .Q_N(\i_ibex/id_stage_i/_0618_ ),
    .Q(\i_ibex/imd_val_q_ex [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[18]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0010_ ),
    .Q_N(\i_ibex/id_stage_i/_0617_ ),
    .Q(\i_ibex/imd_val_q_ex [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[19]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0011_ ),
    .Q_N(\i_ibex/id_stage_i/_0616_ ),
    .Q(\i_ibex/imd_val_q_ex [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[1]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0012_ ),
    .Q_N(\i_ibex/id_stage_i/_0615_ ),
    .Q(\i_ibex/imd_val_q_ex [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[20]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0013_ ),
    .Q_N(\i_ibex/id_stage_i/_0614_ ),
    .Q(\i_ibex/imd_val_q_ex [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[21]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0014_ ),
    .Q_N(\i_ibex/id_stage_i/_0613_ ),
    .Q(\i_ibex/imd_val_q_ex [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[22]_reg  (.CLK(clknet_leaf_0_clk_i_regs),
    .RESET_B(net1553),
    .D(\i_ibex/id_stage_i/_0015_ ),
    .Q_N(\i_ibex/id_stage_i/_0612_ ),
    .Q(\i_ibex/imd_val_q_ex [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[23]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0016_ ),
    .Q_N(\i_ibex/id_stage_i/_0611_ ),
    .Q(\i_ibex/imd_val_q_ex [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[24]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0017_ ),
    .Q_N(\i_ibex/id_stage_i/_0610_ ),
    .Q(\i_ibex/imd_val_q_ex [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[25]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0018_ ),
    .Q_N(\i_ibex/id_stage_i/_0609_ ),
    .Q(\i_ibex/imd_val_q_ex [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[26]_reg  (.CLK(clknet_leaf_0_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0019_ ),
    .Q_N(\i_ibex/id_stage_i/_0608_ ),
    .Q(\i_ibex/imd_val_q_ex [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[27]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0020_ ),
    .Q_N(\i_ibex/id_stage_i/_0607_ ),
    .Q(\i_ibex/imd_val_q_ex [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[28]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0021_ ),
    .Q_N(\i_ibex/id_stage_i/_0606_ ),
    .Q(\i_ibex/imd_val_q_ex [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[29]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0022_ ),
    .Q_N(\i_ibex/id_stage_i/_0605_ ),
    .Q(\i_ibex/imd_val_q_ex [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[2]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0023_ ),
    .Q_N(\i_ibex/id_stage_i/_0604_ ),
    .Q(\i_ibex/imd_val_q_ex [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[30]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0024_ ),
    .Q_N(\i_ibex/id_stage_i/_0603_ ),
    .Q(\i_ibex/imd_val_q_ex [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[31]_reg  (.CLK(clknet_leaf_0_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0025_ ),
    .Q_N(\i_ibex/id_stage_i/_0602_ ),
    .Q(\i_ibex/imd_val_q_ex [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[32]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0026_ ),
    .Q_N(\i_ibex/id_stage_i/_0601_ ),
    .Q(\i_ibex/imd_val_q_ex [32]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[33]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0027_ ),
    .Q_N(\i_ibex/id_stage_i/_0600_ ),
    .Q(\i_ibex/imd_val_q_ex [33]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[34]_reg  (.CLK(clknet_leaf_160_clk_i_regs),
    .RESET_B(net1557),
    .D(\i_ibex/id_stage_i/_0028_ ),
    .Q_N(\i_ibex/id_stage_i/_0599_ ),
    .Q(\i_ibex/imd_val_q_ex [34]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[35]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0029_ ),
    .Q_N(\i_ibex/id_stage_i/_0598_ ),
    .Q(\i_ibex/imd_val_q_ex [35]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[36]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0030_ ),
    .Q_N(\i_ibex/id_stage_i/_0597_ ),
    .Q(\i_ibex/imd_val_q_ex [36]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[37]_reg  (.CLK(clknet_leaf_160_clk_i_regs),
    .RESET_B(net1557),
    .D(\i_ibex/id_stage_i/_0031_ ),
    .Q_N(\i_ibex/id_stage_i/_0596_ ),
    .Q(\i_ibex/imd_val_q_ex [37]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[38]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1556),
    .D(\i_ibex/id_stage_i/_0032_ ),
    .Q_N(\i_ibex/id_stage_i/_0595_ ),
    .Q(\i_ibex/imd_val_q_ex [38]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[39]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0033_ ),
    .Q_N(\i_ibex/id_stage_i/_0594_ ),
    .Q(\i_ibex/imd_val_q_ex [39]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[3]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0034_ ),
    .Q_N(\i_ibex/id_stage_i/_0593_ ),
    .Q(\i_ibex/imd_val_q_ex [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[40]_reg  (.CLK(clknet_leaf_144_clk_i_regs),
    .RESET_B(net1559),
    .D(\i_ibex/id_stage_i/_0035_ ),
    .Q_N(\i_ibex/id_stage_i/_0592_ ),
    .Q(\i_ibex/imd_val_q_ex [40]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[41]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0036_ ),
    .Q_N(\i_ibex/id_stage_i/_0591_ ),
    .Q(\i_ibex/imd_val_q_ex [41]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[42]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0037_ ),
    .Q_N(\i_ibex/id_stage_i/_0590_ ),
    .Q(\i_ibex/imd_val_q_ex [42]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[43]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0038_ ),
    .Q_N(\i_ibex/id_stage_i/_0589_ ),
    .Q(\i_ibex/imd_val_q_ex [43]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[44]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1559),
    .D(\i_ibex/id_stage_i/_0039_ ),
    .Q_N(\i_ibex/id_stage_i/_0588_ ),
    .Q(\i_ibex/imd_val_q_ex [44]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[45]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0040_ ),
    .Q_N(\i_ibex/id_stage_i/_0587_ ),
    .Q(\i_ibex/imd_val_q_ex [45]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[46]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0041_ ),
    .Q_N(\i_ibex/id_stage_i/_0586_ ),
    .Q(\i_ibex/imd_val_q_ex [46]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[47]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0042_ ),
    .Q_N(\i_ibex/id_stage_i/_0585_ ),
    .Q(\i_ibex/imd_val_q_ex [47]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[48]_reg  (.CLK(clknet_leaf_160_clk_i_regs),
    .RESET_B(net1557),
    .D(\i_ibex/id_stage_i/_0043_ ),
    .Q_N(\i_ibex/id_stage_i/_0584_ ),
    .Q(\i_ibex/imd_val_q_ex [48]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[49]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0044_ ),
    .Q_N(\i_ibex/id_stage_i/_0583_ ),
    .Q(\i_ibex/imd_val_q_ex [49]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[4]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0045_ ),
    .Q_N(\i_ibex/id_stage_i/_0582_ ),
    .Q(\i_ibex/imd_val_q_ex [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[50]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0046_ ),
    .Q_N(\i_ibex/id_stage_i/_0581_ ),
    .Q(\i_ibex/imd_val_q_ex [50]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[51]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0047_ ),
    .Q_N(\i_ibex/id_stage_i/_0580_ ),
    .Q(\i_ibex/imd_val_q_ex [51]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[52]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0048_ ),
    .Q_N(\i_ibex/id_stage_i/_0579_ ),
    .Q(\i_ibex/imd_val_q_ex [52]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[53]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0049_ ),
    .Q_N(\i_ibex/id_stage_i/_0578_ ),
    .Q(\i_ibex/imd_val_q_ex [53]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[54]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1556),
    .D(\i_ibex/id_stage_i/_0050_ ),
    .Q_N(\i_ibex/id_stage_i/_0577_ ),
    .Q(\i_ibex/imd_val_q_ex [54]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[55]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0051_ ),
    .Q_N(\i_ibex/id_stage_i/_0576_ ),
    .Q(\i_ibex/imd_val_q_ex [55]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[56]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1557),
    .D(\i_ibex/id_stage_i/_0052_ ),
    .Q_N(\i_ibex/id_stage_i/_0575_ ),
    .Q(\i_ibex/imd_val_q_ex [56]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[57]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0053_ ),
    .Q_N(\i_ibex/id_stage_i/_0574_ ),
    .Q(\i_ibex/imd_val_q_ex [57]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[58]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0054_ ),
    .Q_N(\i_ibex/id_stage_i/_0573_ ),
    .Q(\i_ibex/imd_val_q_ex [58]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[59]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1559),
    .D(\i_ibex/id_stage_i/_0055_ ),
    .Q_N(\i_ibex/id_stage_i/_0572_ ),
    .Q(\i_ibex/imd_val_q_ex [59]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[5]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1527),
    .D(\i_ibex/id_stage_i/_0056_ ),
    .Q_N(\i_ibex/id_stage_i/_0571_ ),
    .Q(\i_ibex/imd_val_q_ex [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[60]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1555),
    .D(\i_ibex/id_stage_i/_0057_ ),
    .Q_N(\i_ibex/id_stage_i/_0570_ ),
    .Q(\i_ibex/imd_val_q_ex [60]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[61]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1558),
    .D(\i_ibex/id_stage_i/_0058_ ),
    .Q_N(\i_ibex/id_stage_i/_0569_ ),
    .Q(\i_ibex/imd_val_q_ex [61]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[62]_reg  (.CLK(clknet_leaf_145_clk_i_regs),
    .RESET_B(net1559),
    .D(\i_ibex/id_stage_i/_0059_ ),
    .Q_N(\i_ibex/id_stage_i/_0568_ ),
    .Q(\i_ibex/imd_val_q_ex [62]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[63]_reg  (.CLK(clknet_leaf_157_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0060_ ),
    .Q_N(\i_ibex/id_stage_i/_0567_ ),
    .Q(\i_ibex/imd_val_q_ex [63]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[64]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0061_ ),
    .Q_N(\i_ibex/id_stage_i/_0566_ ),
    .Q(\i_ibex/imd_val_q_ex [64]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[65]_reg  (.CLK(clknet_leaf_160_clk_i_regs),
    .RESET_B(net1556),
    .D(\i_ibex/id_stage_i/_0062_ ),
    .Q_N(\i_ibex/id_stage_i/_0565_ ),
    .Q(\i_ibex/imd_val_q_ex [65]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[66]_reg  (.CLK(clknet_leaf_158_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0063_ ),
    .Q_N(\i_ibex/id_stage_i/_0564_ ),
    .Q(\i_ibex/imd_val_q_ex [66]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[67]_reg  (.CLK(clknet_leaf_159_clk_i_regs),
    .RESET_B(net1554),
    .D(\i_ibex/id_stage_i/_0064_ ),
    .Q_N(\i_ibex/id_stage_i/_0563_ ),
    .Q(\i_ibex/imd_val_q_ex [67]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[6]_reg  (.CLK(clknet_leaf_161_clk_i_regs),
    .RESET_B(net1523),
    .D(\i_ibex/id_stage_i/_0065_ ),
    .Q_N(\i_ibex/id_stage_i/_0562_ ),
    .Q(\i_ibex/imd_val_q_ex [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[7]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1525),
    .D(\i_ibex/id_stage_i/_0066_ ),
    .Q_N(\i_ibex/id_stage_i/_0561_ ),
    .Q(\i_ibex/imd_val_q_ex [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[8]_reg  (.CLK(clknet_leaf_163_clk_i_regs),
    .RESET_B(net1524),
    .D(\i_ibex/id_stage_i/_0067_ ),
    .Q_N(\i_ibex/id_stage_i/_0560_ ),
    .Q(\i_ibex/imd_val_q_ex [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/id_stage_i/imd_val_q_ex_o[9]_reg  (.CLK(clknet_leaf_162_clk_i_regs),
    .RESET_B(net1526),
    .D(\i_ibex/id_stage_i/_0068_ ),
    .Q_N(\i_ibex/id_stage_i/_0559_ ),
    .Q(\i_ibex/imd_val_q_ex [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/_442_  (.A(\i_ibex/if_stage_i/fetch_err ),
    .B_N(\i_ibex/if_stage_i/fetch_valid ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i_valid_i ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_443_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_084_ ),
    .A(net1122),
    .VSS(VSS));
 sg13g2_buf_2 fanout583 (.A(net585),
    .X(net583),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout582 (.A(\i_ibex/alu_operand_a_ex [30]),
    .X(net582),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout580 (.A(\i_ibex/alu_operand_a_ex [21]),
    .X(net580),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout578 (.A(\i_ibex/alu_operand_a_ex [20]),
    .X(net578),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/if_stage_i/_450_  (.A(\i_ibex/if_stage_i/_084_ ),
    .B(\i_ibex/pc_mux_id [2]),
    .C(\i_ibex/pc_mux_id [0]),
    .D(net1314),
    .Y(\i_ibex/csr_mtvec_init ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_451_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_091_ ),
    .A(net1771),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/_452_  (.A(net623),
    .B(net1307),
    .Y(\i_ibex/if_stage_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/_453_  (.B(\i_ibex/if_stage_i/_092_ ),
    .A(net627),
    .X(\i_ibex/if_stage_i/_093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout576 (.A(\i_ibex/alu_operand_a_ex [19]),
    .X(net576),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_456_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_096_ ),
    .A(net623),
    .VSS(VSS));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/if_stage_i/_458_  (.Y(\i_ibex/if_stage_i/_098_ ),
    .B(net630),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1309));
 sg13g2_buf_2 fanout574 (.A(\i_ibex/alu_operand_a_ex [18]),
    .X(net574),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/if_stage_i/_460_  (.Y(\i_ibex/if_stage_i/_100_ ),
    .B(net1313),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net627));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_462_  (.B1(net1230),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_102_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [31]),
    .A2(net1234));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(\i_ibex/alu_operand_a_ex [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_464_  (.Y(\i_ibex/if_stage_i/_104_ ),
    .B(net1314),
    .A_N(\i_ibex/csr_mepc [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_465_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [32]),
    .A2(\i_ibex/if_stage_i/_104_ ),
    .Y(\i_ibex/if_stage_i/_105_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_466_  (.A2(\i_ibex/if_stage_i/_102_ ),
    .A1(net1239),
    .B1(\i_ibex/if_stage_i/_105_ ),
    .X(\i_ibex/if_stage_i/_106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_467_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_107_ ),
    .A(\i_ibex/csr_mtvec [31]),
    .VSS(VSS));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(\i_ibex/alu_operand_a_ex [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_470_  (.B1(net1314),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_110_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_107_ ),
    .A2(net1342));
 sg13g2_nor2_1 \i_ibex/if_stage_i/_471_  (.A(net630),
    .B(net623),
    .Y(\i_ibex/if_stage_i/_111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/_472_  (.A(net623),
    .B(net1314),
    .X(\i_ibex/if_stage_i/_112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout569 (.A(\i_ibex/alu_operand_a_ex [15]),
    .X(net569),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_474_  (.Y(\i_ibex/if_stage_i/_114_ ),
    .B1(net1221),
    .B2(\i_ibex/csr_mepc [31]),
    .A2(net1226),
    .A1(\i_ibex/if_stage_i/_110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_475_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [31]),
    .B1(\i_ibex/if_stage_i/_106_ ),
    .B2(\i_ibex/if_stage_i/_114_ ),
    .A2(net1187),
    .A1(\i_ibex/if_stage_i/_091_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_476_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_115_ ),
    .A(net1765),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_477_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_116_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [30]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_478_  (.Y(\i_ibex/if_stage_i/_117_ ),
    .B(net1312),
    .A_N(\i_ibex/csr_mepc [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_479_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1520),
    .A2(\i_ibex/if_stage_i/_117_ ),
    .Y(\i_ibex/if_stage_i/_118_ ),
    .B1(net627));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_480_  (.A2(\i_ibex/if_stage_i/_116_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_118_ ),
    .X(\i_ibex/if_stage_i/_119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_481_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_120_ ),
    .A(\i_ibex/csr_mtvec [30]),
    .VSS(VSS));
 sg13g2_buf_2 fanout568 (.A(\i_ibex/alu_operand_a_ex [14]),
    .X(net568),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_483_  (.B1(net1311),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_122_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_120_ ),
    .A2(net1341));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_485_  (.Y(\i_ibex/if_stage_i/_124_ ),
    .B1(\i_ibex/if_stage_i/_122_ ),
    .B2(net1224),
    .A2(net1220),
    .A1(\i_ibex/csr_mepc [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_486_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [30]),
    .B1(\i_ibex/if_stage_i/_119_ ),
    .B2(\i_ibex/if_stage_i/_124_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_487_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_125_ ),
    .A(net1775),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_488_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_126_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [21]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_489_  (.Y(\i_ibex/if_stage_i/_127_ ),
    .B(net1312),
    .A_N(\i_ibex/csr_mepc [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_490_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [22]),
    .A2(\i_ibex/if_stage_i/_127_ ),
    .Y(\i_ibex/if_stage_i/_128_ ),
    .B1(net627));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_491_  (.A2(\i_ibex/if_stage_i/_126_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_128_ ),
    .X(\i_ibex/if_stage_i/_129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_492_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_130_ ),
    .A(\i_ibex/csr_mtvec [21]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_493_  (.B1(net1311),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_131_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_130_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_494_  (.Y(\i_ibex/if_stage_i/_132_ ),
    .B1(\i_ibex/if_stage_i/_131_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_495_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [21]),
    .B1(\i_ibex/if_stage_i/_129_ ),
    .B2(\i_ibex/if_stage_i/_132_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_496_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_133_ ),
    .A(net1762),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_497_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_134_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [20]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_498_  (.Y(\i_ibex/if_stage_i/_135_ ),
    .B(net1312),
    .A_N(\i_ibex/csr_mepc [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_499_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [21]),
    .A2(\i_ibex/if_stage_i/_135_ ),
    .Y(\i_ibex/if_stage_i/_136_ ),
    .B1(net627));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_500_  (.A2(\i_ibex/if_stage_i/_134_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_136_ ),
    .X(\i_ibex/if_stage_i/_137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_501_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_138_ ),
    .A(\i_ibex/csr_mtvec [20]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_502_  (.B1(net1310),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_139_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_138_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_503_  (.Y(\i_ibex/if_stage_i/_140_ ),
    .B1(\i_ibex/if_stage_i/_139_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_504_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [20]),
    .B1(\i_ibex/if_stage_i/_137_ ),
    .B2(\i_ibex/if_stage_i/_140_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_505_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_141_ ),
    .A(net1778),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_506_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_142_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [19]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_507_  (.Y(\i_ibex/if_stage_i/_143_ ),
    .B(net1312),
    .A_N(\i_ibex/csr_mepc [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_508_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [20]),
    .A2(\i_ibex/if_stage_i/_143_ ),
    .Y(\i_ibex/if_stage_i/_144_ ),
    .B1(net627));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_509_  (.A2(\i_ibex/if_stage_i/_142_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_144_ ),
    .X(\i_ibex/if_stage_i/_145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_510_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_146_ ),
    .A(\i_ibex/csr_mtvec [19]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_511_  (.B1(net1310),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_147_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_146_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_512_  (.Y(\i_ibex/if_stage_i/_148_ ),
    .B1(\i_ibex/if_stage_i/_147_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_513_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [19]),
    .B1(\i_ibex/if_stage_i/_145_ ),
    .B2(\i_ibex/if_stage_i/_148_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_514_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_149_ ),
    .A(net1760),
    .VSS(VSS));
 sg13g2_buf_2 fanout566 (.A(\i_ibex/alu_operand_a_ex [13]),
    .X(net566),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_516_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_151_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [18]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_517_  (.Y(\i_ibex/if_stage_i/_152_ ),
    .B(net1311),
    .A_N(\i_ibex/csr_mepc [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout565 (.A(net566),
    .X(net565),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_519_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [19]),
    .A2(\i_ibex/if_stage_i/_152_ ),
    .Y(\i_ibex/if_stage_i/_154_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_520_  (.A2(\i_ibex/if_stage_i/_151_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_154_ ),
    .X(\i_ibex/if_stage_i/_155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_521_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_156_ ),
    .A(\i_ibex/csr_mtvec [18]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_522_  (.B1(net1310),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_157_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_156_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_523_  (.Y(\i_ibex/if_stage_i/_158_ ),
    .B1(\i_ibex/if_stage_i/_157_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_524_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [18]),
    .B1(\i_ibex/if_stage_i/_155_ ),
    .B2(\i_ibex/if_stage_i/_158_ ),
    .A2(net1186),
    .A1(\i_ibex/if_stage_i/_149_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_525_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_159_ ),
    .A(net1773),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_526_  (.B1(net1230),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_160_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [17]),
    .A2(net1234));
 sg13g2_buf_2 fanout564 (.A(\i_ibex/alu_operand_a_ex [12]),
    .X(net564),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_528_  (.Y(\i_ibex/if_stage_i/_162_ ),
    .B(net1315),
    .A_N(\i_ibex/csr_mepc [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_529_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [18]),
    .A2(\i_ibex/if_stage_i/_162_ ),
    .Y(\i_ibex/if_stage_i/_163_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_530_  (.A2(\i_ibex/if_stage_i/_160_ ),
    .A1(net1239),
    .B1(\i_ibex/if_stage_i/_163_ ),
    .X(\i_ibex/if_stage_i/_164_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_531_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_165_ ),
    .A(\i_ibex/csr_mtvec [17]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_532_  (.B1(net1314),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_166_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_165_ ),
    .A2(net1342));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_533_  (.Y(\i_ibex/if_stage_i/_167_ ),
    .B1(\i_ibex/if_stage_i/_166_ ),
    .B2(net1226),
    .A2(net1221),
    .A1(\i_ibex/csr_mepc [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_534_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [17]),
    .B1(\i_ibex/if_stage_i/_164_ ),
    .B2(\i_ibex/if_stage_i/_167_ ),
    .A2(net1187),
    .A1(\i_ibex/if_stage_i/_159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_535_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_168_ ),
    .A(net1782),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_536_  (.B1(net1229),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_169_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [16]),
    .A2(net1233));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_537_  (.Y(\i_ibex/if_stage_i/_170_ ),
    .B(net1313),
    .A_N(\i_ibex/csr_mepc [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_538_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [17]),
    .A2(\i_ibex/if_stage_i/_170_ ),
    .Y(\i_ibex/if_stage_i/_171_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_539_  (.A2(\i_ibex/if_stage_i/_169_ ),
    .A1(net1238),
    .B1(\i_ibex/if_stage_i/_171_ ),
    .X(\i_ibex/if_stage_i/_172_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_540_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_173_ ),
    .A(\i_ibex/csr_mtvec [16]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_541_  (.B1(net1313),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_174_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_173_ ),
    .A2(net1341));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_542_  (.Y(\i_ibex/if_stage_i/_175_ ),
    .B1(\i_ibex/if_stage_i/_174_ ),
    .B2(net1225),
    .A2(net1220),
    .A1(\i_ibex/csr_mepc [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_543_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [16]),
    .B1(\i_ibex/if_stage_i/_172_ ),
    .B2(\i_ibex/if_stage_i/_175_ ),
    .A2(net1186),
    .A1(\i_ibex/if_stage_i/_168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_544_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_176_ ),
    .A(net1780),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_545_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_177_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [15]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_546_  (.Y(\i_ibex/if_stage_i/_178_ ),
    .B(net1307),
    .A_N(\i_ibex/csr_mepc [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_547_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [16]),
    .A2(\i_ibex/if_stage_i/_178_ ),
    .Y(\i_ibex/if_stage_i/_179_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_548_  (.A2(\i_ibex/if_stage_i/_177_ ),
    .A1(net1236),
    .B1(\i_ibex/if_stage_i/_179_ ),
    .X(\i_ibex/if_stage_i/_180_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_549_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_181_ ),
    .A(\i_ibex/csr_mtvec [15]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_550_  (.B1(net1314),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_182_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_181_ ),
    .A2(net1339));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_551_  (.Y(\i_ibex/if_stage_i/_183_ ),
    .B1(\i_ibex/if_stage_i/_182_ ),
    .B2(net1223),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_552_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [15]),
    .B1(\i_ibex/if_stage_i/_180_ ),
    .B2(\i_ibex/if_stage_i/_183_ ),
    .A2(net1184),
    .A1(\i_ibex/if_stage_i/_176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_553_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_184_ ),
    .A(boot_addr_i[14]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_554_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_185_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [14]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_555_  (.Y(\i_ibex/if_stage_i/_186_ ),
    .B(net1307),
    .A_N(\i_ibex/csr_mepc [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_556_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [15]),
    .A2(\i_ibex/if_stage_i/_186_ ),
    .Y(\i_ibex/if_stage_i/_187_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_557_  (.A2(\i_ibex/if_stage_i/_185_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_187_ ),
    .X(\i_ibex/if_stage_i/_188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_558_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_189_ ),
    .A(\i_ibex/csr_mtvec [14]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_559_  (.B1(net1305),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_190_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_189_ ),
    .A2(net1338));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_560_  (.Y(\i_ibex/if_stage_i/_191_ ),
    .B1(\i_ibex/if_stage_i/_190_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_561_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [14]),
    .B1(\i_ibex/if_stage_i/_188_ ),
    .B2(\i_ibex/if_stage_i/_191_ ),
    .A2(net1182),
    .A1(\i_ibex/if_stage_i/_184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_562_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_192_ ),
    .A(net1774),
    .VSS(VSS));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout561 (.A(\i_ibex/alu_operand_a_ex [29]),
    .X(net561),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_566_  (.B1(\i_ibex/if_stage_i/_100_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_196_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [13]),
    .A2(\i_ibex/if_stage_i/_098_ ));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_567_  (.Y(\i_ibex/if_stage_i/_197_ ),
    .B(net1307),
    .A_N(\i_ibex/csr_mepc [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_568_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [14]),
    .A2(\i_ibex/if_stage_i/_197_ ),
    .Y(\i_ibex/if_stage_i/_198_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_569_  (.A2(\i_ibex/if_stage_i/_196_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_198_ ),
    .X(\i_ibex/if_stage_i/_199_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_571_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_201_ ),
    .A(\i_ibex/csr_mtvec [13]),
    .VSS(VSS));
 sg13g2_buf_2 fanout559 (.A(\i_ibex/alu_operand_a_ex [11]),
    .X(net559),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_573_  (.B1(net1308),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_203_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_201_ ),
    .A2(net1338));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_574_  (.Y(\i_ibex/if_stage_i/_204_ ),
    .B1(\i_ibex/if_stage_i/_203_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_575_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [13]),
    .B1(\i_ibex/if_stage_i/_199_ ),
    .B2(\i_ibex/if_stage_i/_204_ ),
    .A2(net1183),
    .A1(\i_ibex/if_stage_i/_192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_576_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_205_ ),
    .A(boot_addr_i[12]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_577_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_206_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [12]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_578_  (.Y(\i_ibex/if_stage_i/_207_ ),
    .B(net1306),
    .A_N(\i_ibex/csr_mepc [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_579_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [13]),
    .A2(\i_ibex/if_stage_i/_207_ ),
    .Y(\i_ibex/if_stage_i/_208_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_580_  (.A2(\i_ibex/if_stage_i/_206_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_208_ ),
    .X(\i_ibex/if_stage_i/_209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_581_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_210_ ),
    .A(\i_ibex/csr_mtvec [12]),
    .VSS(VSS));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_583_  (.B1(net1306),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_212_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_210_ ),
    .A2(net1339));
 sg13g2_buf_1 fanout557 (.A(\i_ibex/alu_operand_a_ex [10]),
    .X(net557),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_585_  (.Y(\i_ibex/if_stage_i/_214_ ),
    .B1(\i_ibex/if_stage_i/_212_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_586_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [12]),
    .B1(\i_ibex/if_stage_i/_209_ ),
    .B2(\i_ibex/if_stage_i/_214_ ),
    .A2(net1182),
    .A1(\i_ibex/if_stage_i/_205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_587_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_215_ ),
    .A(net1776),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_588_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_216_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [29]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_589_  (.Y(\i_ibex/if_stage_i/_217_ ),
    .B(net1308),
    .A_N(\i_ibex/csr_mepc [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_590_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1518),
    .A2(\i_ibex/if_stage_i/_217_ ),
    .Y(\i_ibex/if_stage_i/_218_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_591_  (.A2(\i_ibex/if_stage_i/_216_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_218_ ),
    .X(\i_ibex/if_stage_i/_219_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_592_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_220_ ),
    .A(\i_ibex/csr_mtvec [29]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_593_  (.B1(net1308),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_221_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_220_ ),
    .A2(net1338));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_594_  (.Y(\i_ibex/if_stage_i/_222_ ),
    .B1(\i_ibex/if_stage_i/_221_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_595_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [29]),
    .B1(\i_ibex/if_stage_i/_219_ ),
    .B2(\i_ibex/if_stage_i/_222_ ),
    .A2(net1183),
    .A1(\i_ibex/if_stage_i/_215_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_596_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_223_ ),
    .A(net1763),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_597_  (.Y(\i_ibex/if_stage_i/_224_ ),
    .A(\i_ibex/csr_mepc [11]),
    .B(net1307),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/_598_  (.A(net623),
    .B_N(net1307),
    .Y(\i_ibex/if_stage_i/_225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_599_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net623),
    .A2(\i_ibex/if_stage_i/_224_ ),
    .Y(\i_ibex/if_stage_i/_226_ ),
    .B1(\i_ibex/if_stage_i/_225_ ));
 sg13g2_nand3b_1 \i_ibex/if_stage_i/_600_  (.B(net630),
    .C(\i_ibex/if_stage_i/_092_ ),
    .Y(\i_ibex/if_stage_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/csr_depc [11]));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_601_  (.B1(\i_ibex/if_stage_i/_227_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_228_ ),
    .VSS(VSS),
    .A1(net627),
    .A2(\i_ibex/if_stage_i/_226_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_602_  (.B1(\i_ibex/if_stage_i/_225_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_229_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_mtvec [11]),
    .A2(net1338));
 sg13g2_nand3b_1 \i_ibex/if_stage_i/_603_  (.B(net623),
    .C(\i_ibex/ex_block_i/alu_adder_result_ext [12]),
    .Y(\i_ibex/if_stage_i/_230_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1307));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_604_  (.A2(\i_ibex/if_stage_i/_230_ ),
    .A1(\i_ibex/if_stage_i/_229_ ),
    .B1(net630),
    .X(\i_ibex/if_stage_i/_231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_605_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [11]),
    .B1(\i_ibex/if_stage_i/_228_ ),
    .B2(\i_ibex/if_stage_i/_231_ ),
    .A2(net1182),
    .A1(\i_ibex/if_stage_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_606_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_232_ ),
    .A(boot_addr_i[10]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_607_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_233_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [10]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_608_  (.Y(\i_ibex/if_stage_i/_234_ ),
    .B(net1306),
    .A_N(\i_ibex/csr_mepc [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_609_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [11]),
    .A2(\i_ibex/if_stage_i/_234_ ),
    .Y(\i_ibex/if_stage_i/_235_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_610_  (.A2(\i_ibex/if_stage_i/_233_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_235_ ),
    .X(\i_ibex/if_stage_i/_236_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_611_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_237_ ),
    .A(\i_ibex/csr_mtvec [10]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_612_  (.B1(net1306),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_238_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_237_ ),
    .A2(net1339));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_613_  (.Y(\i_ibex/if_stage_i/_239_ ),
    .B1(\i_ibex/if_stage_i/_238_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_614_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .B1(\i_ibex/if_stage_i/_236_ ),
    .B2(\i_ibex/if_stage_i/_239_ ),
    .A2(net1183),
    .A1(\i_ibex/if_stage_i/_232_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_615_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_240_ ),
    .A(net1761),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_616_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_241_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [9]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_617_  (.Y(\i_ibex/if_stage_i/_242_ ),
    .B(net1306),
    .A_N(\i_ibex/csr_mepc [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_618_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [10]),
    .A2(\i_ibex/if_stage_i/_242_ ),
    .Y(\i_ibex/if_stage_i/_243_ ),
    .B1(net628));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_619_  (.A2(\i_ibex/if_stage_i/_241_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_243_ ),
    .X(\i_ibex/if_stage_i/_244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_620_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_245_ ),
    .A(\i_ibex/csr_mtvec [9]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_621_  (.B1(net1306),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_246_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_245_ ),
    .A2(net1338));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_622_  (.Y(\i_ibex/if_stage_i/_247_ ),
    .B1(\i_ibex/if_stage_i/_246_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_623_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [9]),
    .B1(\i_ibex/if_stage_i/_244_ ),
    .B2(\i_ibex/if_stage_i/_247_ ),
    .A2(net1183),
    .A1(\i_ibex/if_stage_i/_240_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_624_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_248_ ),
    .A(net1779),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_625_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_249_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [8]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_626_  (.Y(\i_ibex/if_stage_i/_250_ ),
    .B(net1308),
    .A_N(\i_ibex/csr_mepc [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_628_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [9]),
    .A2(\i_ibex/if_stage_i/_250_ ),
    .Y(\i_ibex/if_stage_i/_252_ ),
    .B1(net630));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_629_  (.A2(\i_ibex/if_stage_i/_249_ ),
    .A1(net1235),
    .B1(\i_ibex/if_stage_i/_252_ ),
    .X(\i_ibex/if_stage_i/_253_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_630_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_254_ ),
    .A(\i_ibex/csr_mtvec [8]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_631_  (.B1(net1308),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_255_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_254_ ),
    .A2(net1338));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_632_  (.Y(\i_ibex/if_stage_i/_256_ ),
    .B1(\i_ibex/if_stage_i/_255_ ),
    .B2(net1222),
    .A2(net1218),
    .A1(\i_ibex/csr_mepc [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_633_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [8]),
    .B1(\i_ibex/if_stage_i/_253_ ),
    .B2(\i_ibex/if_stage_i/_256_ ),
    .A2(net1183),
    .A1(\i_ibex/if_stage_i/_248_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_634_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_257_ ),
    .A(net1338),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/if_stage_i/_635_  (.A(net1307),
    .B(\i_ibex/exc_pc_mux_id [0]),
    .C(\i_ibex/if_stage_i/_257_ ),
    .D(net1222),
    .X(\i_ibex/if_stage_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_636_  (.Y(\i_ibex/if_stage_i/_259_ ),
    .A(\i_ibex/exc_cause [5]),
    .B(\i_ibex/if_stage_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/if_stage_i/_637_  (.A(net630),
    .B(\i_ibex/if_stage_i/_092_ ),
    .X(\i_ibex/if_stage_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_638_  (.A0(\i_ibex/ex_block_i/alu_adder_result_ext [8]),
    .A1(\i_ibex/csr_mepc [7]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/if_stage_i/_639_  (.A(\i_ibex/pc_mux_id [2]),
    .B(net1235),
    .Y(\i_ibex/if_stage_i/_262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_640_  (.Y(\i_ibex/if_stage_i/_263_ ),
    .B1(\i_ibex/if_stage_i/_261_ ),
    .B2(\i_ibex/if_stage_i/_262_ ),
    .A2(\i_ibex/if_stage_i/_260_ ),
    .A1(\i_ibex/csr_depc [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/_641_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1182),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [7]),
    .A2(\i_ibex/if_stage_i/_263_ ),
    .A1(\i_ibex/if_stage_i/_259_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_642_  (.Y(\i_ibex/if_stage_i/_264_ ),
    .A(\i_ibex/exc_cause [4]),
    .B(\i_ibex/if_stage_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_643_  (.A0(\i_ibex/ex_block_i/alu_adder_result_ext [7]),
    .A1(\i_ibex/csr_mepc [6]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_265_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_644_  (.Y(\i_ibex/if_stage_i/_266_ ),
    .B1(\i_ibex/if_stage_i/_262_ ),
    .B2(\i_ibex/if_stage_i/_265_ ),
    .A2(\i_ibex/if_stage_i/_260_ ),
    .A1(\i_ibex/csr_depc [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/_645_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1182),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [6]),
    .A2(\i_ibex/if_stage_i/_266_ ),
    .A1(\i_ibex/if_stage_i/_264_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_646_  (.Y(\i_ibex/if_stage_i/_267_ ),
    .A(\i_ibex/exc_cause [3]),
    .B(\i_ibex/if_stage_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_647_  (.A0(\i_ibex/ex_block_i/alu_adder_result_ext [6]),
    .A1(\i_ibex/csr_mepc [5]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_648_  (.Y(\i_ibex/if_stage_i/_269_ ),
    .B1(\i_ibex/if_stage_i/_262_ ),
    .B2(\i_ibex/if_stage_i/_268_ ),
    .A2(\i_ibex/if_stage_i/_260_ ),
    .A1(\i_ibex/csr_depc [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/_649_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1182),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [5]),
    .A2(\i_ibex/if_stage_i/_269_ ),
    .A1(\i_ibex/if_stage_i/_267_ ));
 sg13g2_or2_1 \i_ibex/if_stage_i/_650_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/_270_ ),
    .B(\i_ibex/exc_cause [2]),
    .A(net1338));
 sg13g2_and2_1 \i_ibex/if_stage_i/_651_  (.A(\i_ibex/exc_pc_mux_id [0]),
    .B(\i_ibex/if_stage_i/_225_ ),
    .X(\i_ibex/if_stage_i/_271_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_652_  (.A0(\i_ibex/ex_block_i/alu_adder_result_ext [5]),
    .A1(\i_ibex/csr_mepc [4]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_272_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_653_  (.Y(\i_ibex/if_stage_i/_273_ ),
    .B1(\i_ibex/if_stage_i/_272_ ),
    .B2(net623),
    .A2(\i_ibex/if_stage_i/_271_ ),
    .A1(\i_ibex/if_stage_i/_270_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_654_  (.Y(\i_ibex/if_stage_i/_274_ ),
    .A(\i_ibex/csr_depc [4]),
    .B(\i_ibex/if_stage_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_655_  (.B1(\i_ibex/if_stage_i/_274_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [4]),
    .VSS(VSS),
    .A1(net627),
    .A2(\i_ibex/if_stage_i/_273_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_656_  (.Y(\i_ibex/if_stage_i/_275_ ),
    .A(\i_ibex/exc_cause [1]),
    .B(\i_ibex/if_stage_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_657_  (.A0(\i_ibex/ex_block_i/alu_adder_result_ext [4]),
    .A1(\i_ibex/csr_mepc [3]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_276_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_658_  (.Y(\i_ibex/if_stage_i/_277_ ),
    .B1(\i_ibex/if_stage_i/_262_ ),
    .B2(\i_ibex/if_stage_i/_276_ ),
    .A2(\i_ibex/if_stage_i/_260_ ),
    .A1(\i_ibex/csr_depc [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/_659_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1182),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [3]),
    .A2(\i_ibex/if_stage_i/_277_ ),
    .A1(\i_ibex/if_stage_i/_275_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_660_  (.Y(\i_ibex/if_stage_i/_278_ ),
    .A(\i_ibex/exc_cause [0]),
    .B(\i_ibex/if_stage_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_661_  (.A0(\i_ibex/ex_block_i/alu_adder_result_ext [3]),
    .A1(\i_ibex/csr_mepc [2]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_279_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_662_  (.Y(\i_ibex/if_stage_i/_280_ ),
    .B1(\i_ibex/if_stage_i/_262_ ),
    .B2(\i_ibex/if_stage_i/_279_ ),
    .A2(\i_ibex/if_stage_i/_260_ ),
    .A1(\i_ibex/csr_depc [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/_663_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1182),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [2]),
    .A2(\i_ibex/if_stage_i/_280_ ),
    .A1(\i_ibex/if_stage_i/_278_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/_664_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_281_ ),
    .A(net1777),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_665_  (.B1(net1230),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_282_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [28]),
    .A2(net1234));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_666_  (.Y(\i_ibex/if_stage_i/_283_ ),
    .B(net1314),
    .A_N(\i_ibex/csr_mepc [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_667_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1519),
    .A2(\i_ibex/if_stage_i/_283_ ),
    .Y(\i_ibex/if_stage_i/_284_ ),
    .B1(net630));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_668_  (.A2(\i_ibex/if_stage_i/_282_ ),
    .A1(net1236),
    .B1(\i_ibex/if_stage_i/_284_ ),
    .X(\i_ibex/if_stage_i/_285_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_669_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_286_ ),
    .A(\i_ibex/csr_mtvec [28]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_670_  (.B1(net1314),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_287_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_286_ ),
    .A2(net1339));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_671_  (.Y(\i_ibex/if_stage_i/_288_ ),
    .B1(\i_ibex/if_stage_i/_287_ ),
    .B2(net1223),
    .A2(net1221),
    .A1(\i_ibex/csr_mepc [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_672_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [28]),
    .B1(\i_ibex/if_stage_i/_285_ ),
    .B2(\i_ibex/if_stage_i/_288_ ),
    .A2(net1184),
    .A1(\i_ibex/if_stage_i/_281_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_673_  (.A0(net435),
    .A1(\i_ibex/csr_mepc [1]),
    .S(net1305),
    .X(\i_ibex/if_stage_i/_289_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_674_  (.Y(\i_ibex/if_stage_i/_290_ ),
    .B1(\i_ibex/if_stage_i/_262_ ),
    .B2(\i_ibex/if_stage_i/_289_ ),
    .A2(\i_ibex/if_stage_i/_260_ ),
    .A1(\i_ibex/csr_depc [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_675_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/fetch_addr_n [1]),
    .A(\i_ibex/if_stage_i/_290_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_676_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_291_ ),
    .A(net1781),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_677_  (.B1(net1227),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_292_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [27]),
    .A2(net1231));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_678_  (.Y(\i_ibex/if_stage_i/_293_ ),
    .B(net1309),
    .A_N(\i_ibex/csr_mepc [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_679_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [28]),
    .A2(\i_ibex/if_stage_i/_293_ ),
    .Y(\i_ibex/if_stage_i/_294_ ),
    .B1(net630));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_680_  (.A2(\i_ibex/if_stage_i/_292_ ),
    .A1(net1236),
    .B1(\i_ibex/if_stage_i/_294_ ),
    .X(\i_ibex/if_stage_i/_295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_681_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_296_ ),
    .A(\i_ibex/csr_mtvec [27]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_682_  (.B1(net1309),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_297_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_296_ ),
    .A2(net1342));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_683_  (.Y(\i_ibex/if_stage_i/_298_ ),
    .B1(\i_ibex/if_stage_i/_297_ ),
    .B2(net1223),
    .A2(net1221),
    .A1(\i_ibex/csr_mepc [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_684_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [27]),
    .B1(\i_ibex/if_stage_i/_295_ ),
    .B2(\i_ibex/if_stage_i/_298_ ),
    .A2(net1184),
    .A1(\i_ibex/if_stage_i/_291_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_685_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_299_ ),
    .A(net1770),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_686_  (.B1(net1229),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_300_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [26]),
    .A2(net1233));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_687_  (.Y(\i_ibex/if_stage_i/_301_ ),
    .B(net1310),
    .A_N(\i_ibex/csr_mepc [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_688_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [27]),
    .A2(\i_ibex/if_stage_i/_301_ ),
    .Y(\i_ibex/if_stage_i/_302_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_689_  (.A2(\i_ibex/if_stage_i/_300_ ),
    .A1(net1238),
    .B1(\i_ibex/if_stage_i/_302_ ),
    .X(\i_ibex/if_stage_i/_303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_690_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_304_ ),
    .A(\i_ibex/csr_mtvec [26]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_691_  (.B1(net1311),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_305_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_304_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_692_  (.Y(\i_ibex/if_stage_i/_306_ ),
    .B1(\i_ibex/if_stage_i/_305_ ),
    .B2(net1225),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_693_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [26]),
    .B1(\i_ibex/if_stage_i/_303_ ),
    .B2(\i_ibex/if_stage_i/_306_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_299_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_694_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_307_ ),
    .A(net1759),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_695_  (.B1(net1229),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_308_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [25]),
    .A2(net1233));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_696_  (.Y(\i_ibex/if_stage_i/_309_ ),
    .B(net1310),
    .A_N(\i_ibex/csr_mepc [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_697_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [26]),
    .A2(\i_ibex/if_stage_i/_309_ ),
    .Y(\i_ibex/if_stage_i/_310_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_698_  (.A2(\i_ibex/if_stage_i/_308_ ),
    .A1(net1238),
    .B1(\i_ibex/if_stage_i/_310_ ),
    .X(\i_ibex/if_stage_i/_311_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_699_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_312_ ),
    .A(\i_ibex/csr_mtvec [25]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_700_  (.B1(net1310),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_313_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_312_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_701_  (.Y(\i_ibex/if_stage_i/_314_ ),
    .B1(\i_ibex/if_stage_i/_313_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_702_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [25]),
    .B1(\i_ibex/if_stage_i/_311_ ),
    .B2(\i_ibex/if_stage_i/_314_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_307_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_703_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_315_ ),
    .A(net1766),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_704_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_316_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [24]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_705_  (.Y(\i_ibex/if_stage_i/_317_ ),
    .B(net1310),
    .A_N(\i_ibex/csr_mepc [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_706_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [25]),
    .A2(\i_ibex/if_stage_i/_317_ ),
    .Y(\i_ibex/if_stage_i/_318_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_707_  (.A2(\i_ibex/if_stage_i/_316_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_318_ ),
    .X(\i_ibex/if_stage_i/_319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_708_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_320_ ),
    .A(\i_ibex/csr_mtvec [24]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_709_  (.B1(net1310),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_321_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_320_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_710_  (.Y(\i_ibex/if_stage_i/_322_ ),
    .B1(\i_ibex/if_stage_i/_321_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_711_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [24]),
    .B1(\i_ibex/if_stage_i/_319_ ),
    .B2(\i_ibex/if_stage_i/_322_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_712_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_323_ ),
    .A(net1768),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_713_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_324_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [23]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_714_  (.Y(\i_ibex/if_stage_i/_325_ ),
    .B(net1312),
    .A_N(\i_ibex/csr_mepc [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_715_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [24]),
    .A2(\i_ibex/if_stage_i/_325_ ),
    .Y(\i_ibex/if_stage_i/_326_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_716_  (.A2(\i_ibex/if_stage_i/_324_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_326_ ),
    .X(\i_ibex/if_stage_i/_327_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_717_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_328_ ),
    .A(\i_ibex/csr_mtvec [23]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_718_  (.B1(net1312),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_329_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_328_ ),
    .A2(net1340));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_719_  (.Y(\i_ibex/if_stage_i/_330_ ),
    .B1(\i_ibex/if_stage_i/_329_ ),
    .B2(net1224),
    .A2(net1219),
    .A1(\i_ibex/csr_mepc [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_720_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .B1(\i_ibex/if_stage_i/_327_ ),
    .B2(\i_ibex/if_stage_i/_330_ ),
    .A2(net1185),
    .A1(\i_ibex/if_stage_i/_323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_721_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_331_ ),
    .A(net1772),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_722_  (.B1(net1228),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_332_ ),
    .VSS(VSS),
    .A1(\i_ibex/csr_depc [22]),
    .A2(net1232));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_723_  (.Y(\i_ibex/if_stage_i/_333_ ),
    .B(net1312),
    .A_N(\i_ibex/csr_mepc [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/_724_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [23]),
    .A2(\i_ibex/if_stage_i/_333_ ),
    .Y(\i_ibex/if_stage_i/_334_ ),
    .B1(net629));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_725_  (.A2(\i_ibex/if_stage_i/_332_ ),
    .A1(net1237),
    .B1(\i_ibex/if_stage_i/_334_ ),
    .X(\i_ibex/if_stage_i/_335_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/_726_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/_336_ ),
    .A(\i_ibex/csr_mtvec [22]),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_727_  (.B1(net1312),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/_337_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/_336_ ),
    .A2(net1341));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_728_  (.Y(\i_ibex/if_stage_i/_338_ ),
    .B1(\i_ibex/if_stage_i/_337_ ),
    .B2(net1225),
    .A2(net1220),
    .A1(\i_ibex/csr_mepc [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/_729_  (.Y(\i_ibex/if_stage_i/fetch_addr_n [22]),
    .B1(\i_ibex/if_stage_i/_335_ ),
    .B2(\i_ibex/if_stage_i/_338_ ),
    .A2(net1186),
    .A1(\i_ibex/if_stage_i/_331_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/_730_  (.Y(\i_ibex/if_stage_i/_339_ ),
    .A(\i_ibex/if_stage_i/fetch_valid ),
    .B(\i_ibex/id_in_ready ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_8 \i_ibex/if_stage_i/_731_  (.Y(\i_ibex/if_stage_i/_340_ ),
    .A(\i_ibex/if_stage_i/_339_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout555 (.A(\i_ibex/alu_operand_a_ex [9]),
    .X(net555),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_734_  (.A0(\i_ibex/illegal_c_insn_id ),
    .A1(\i_ibex/if_stage_i/illegal_c_insn ),
    .S(net835),
    .X(\i_ibex/if_stage_i/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/if_stage_i/_735_  (.B(\i_ibex/pc_if [2]),
    .C(net42),
    .Y(\i_ibex/if_stage_i/_342_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/if_stage_i/instr_is_compressed ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/_736_  (.A(\i_ibex/if_stage_i/fetch_err ),
    .B(net43),
    .Y(\i_ibex/if_stage_i/_343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/_737_  (.Y(\i_ibex/if_stage_i/_344_ ),
    .A(\i_ibex/if_stage_i/_342_ ),
    .B(\i_ibex/if_stage_i/_343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_738_  (.A0(\i_ibex/instr_fetch_err ),
    .A1(\i_ibex/if_stage_i/_344_ ),
    .S(net837),
    .X(\i_ibex/if_stage_i/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/_739_  (.A(\i_ibex/if_stage_i/fetch_err_plus2 ),
    .B_N(\i_ibex/if_stage_i/_342_ ),
    .Y(\i_ibex/if_stage_i/_345_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/_740_  (.A(net44),
    .B(\i_ibex/if_stage_i/_339_ ),
    .C(\i_ibex/if_stage_i/_345_ ),
    .Y(\i_ibex/if_stage_i/_346_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/_741_  (.A2(\i_ibex/if_stage_i/_339_ ),
    .A1(\i_ibex/instr_fetch_err_plus2 ),
    .B1(\i_ibex/if_stage_i/_346_ ),
    .X(\i_ibex/if_stage_i/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_742_  (.A0(\i_ibex/if_stage_i/instr_is_compressed ),
    .A1(\i_ibex/instr_is_compressed_id ),
    .S(\i_ibex/if_stage_i/_339_ ),
    .X(\i_ibex/if_stage_i/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_743_  (.A0(\i_ibex/instr_rdata_id [0]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [0]),
    .S(net829),
    .X(\i_ibex/if_stage_i/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_744_  (.A0(\i_ibex/id_stage_i/imm_s_type [3]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [10]),
    .S(net829),
    .X(\i_ibex/if_stage_i/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_745_  (.A0(\i_ibex/id_stage_i/imm_s_type [4]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [11]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_746_  (.A0(\i_ibex/id_stage_i/imm_u_type [12]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [12]),
    .S(net831),
    .X(\i_ibex/if_stage_i/_007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_747_  (.A0(\i_ibex/id_stage_i/imm_u_type [13]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [13]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_748_  (.A0(\i_ibex/id_stage_i/imm_u_type [14]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [14]),
    .S(net836),
    .X(\i_ibex/if_stage_i/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_749_  (.A0(\i_ibex/id_stage_i/zimm_rs1_type [0]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [15]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout553 (.A(\i_ibex/alu_operand_a_ex [8]),
    .X(net553),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_751_  (.A0(\i_ibex/id_stage_i/zimm_rs1_type [1]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [16]),
    .S(net829),
    .X(\i_ibex/if_stage_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_752_  (.A0(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [17]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_753_  (.A0(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [18]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_754_  (.A0(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [19]),
    .S(net834),
    .X(\i_ibex/if_stage_i/_014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_755_  (.A0(\i_ibex/instr_rdata_id [1]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [1]),
    .S(net831),
    .X(\i_ibex/if_stage_i/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_756_  (.A0(net762),
    .A1(\i_ibex/if_stage_i/instr_decompressed [20]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_757_  (.A0(net758),
    .A1(\i_ibex/if_stage_i/instr_decompressed [21]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_758_  (.A0(net756),
    .A1(\i_ibex/if_stage_i/instr_decompressed [22]),
    .S(net836),
    .X(\i_ibex/if_stage_i/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_759_  (.A0(\i_ibex/id_stage_i/imm_u_type [23]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [23]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_760_  (.A0(\i_ibex/id_stage_i/imm_u_type [24]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [24]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_762_  (.A0(\i_ibex/id_stage_i/imm_u_type [25]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [25]),
    .S(net831),
    .X(\i_ibex/if_stage_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_763_  (.A0(net749),
    .A1(\i_ibex/if_stage_i/instr_decompressed [26]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_764_  (.A0(\i_ibex/id_stage_i/imm_u_type [27]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [27]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_765_  (.A0(\i_ibex/id_stage_i/imm_u_type [28]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [28]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_766_  (.A0(\i_ibex/id_stage_i/imm_u_type [29]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [29]),
    .S(net832),
    .X(\i_ibex/if_stage_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_767_  (.A0(\i_ibex/instr_rdata_id [2]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [2]),
    .S(net832),
    .X(\i_ibex/if_stage_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_768_  (.A0(\i_ibex/id_stage_i/imm_u_type [30]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [30]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_769_  (.A0(net733),
    .A1(\i_ibex/if_stage_i/instr_decompressed [31]),
    .S(net831),
    .X(\i_ibex/if_stage_i/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_770_  (.A0(\i_ibex/instr_rdata_id [3]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [3]),
    .S(net835),
    .X(\i_ibex/if_stage_i/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_771_  (.A0(net718),
    .A1(\i_ibex/if_stage_i/instr_decompressed [4]),
    .S(net836),
    .X(\i_ibex/if_stage_i/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout551 (.A(\i_ibex/alu_operand_a_ex [7]),
    .X(net551),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_773_  (.A0(\i_ibex/instr_rdata_id [5]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [5]),
    .S(net836),
    .X(\i_ibex/if_stage_i/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_774_  (.A0(net711),
    .A1(\i_ibex/if_stage_i/instr_decompressed [6]),
    .S(net836),
    .X(\i_ibex/if_stage_i/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_775_  (.A0(\i_ibex/id_stage_i/imm_s_type [0]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [7]),
    .S(net829),
    .X(\i_ibex/if_stage_i/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_776_  (.A0(\i_ibex/id_stage_i/imm_s_type [1]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [8]),
    .S(net833),
    .X(\i_ibex/if_stage_i/_034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_777_  (.A0(\i_ibex/id_stage_i/imm_s_type [2]),
    .A1(\i_ibex/if_stage_i/instr_decompressed [9]),
    .S(net829),
    .X(\i_ibex/if_stage_i/_035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_778_  (.A0(\i_ibex/instr_rdata_c_id [0]),
    .A1(net636),
    .S(net829),
    .X(\i_ibex/if_stage_i/_036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_779_  (.A0(\i_ibex/instr_rdata_c_id [10]),
    .A1(net1359),
    .S(net830),
    .X(\i_ibex/if_stage_i/_037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_780_  (.A0(\i_ibex/instr_rdata_c_id [11]),
    .A1(net644),
    .S(net830),
    .X(\i_ibex/if_stage_i/_038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_781_  (.A0(\i_ibex/instr_rdata_c_id [12]),
    .A1(net646),
    .S(net831),
    .X(\i_ibex/if_stage_i/_039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_782_  (.A0(\i_ibex/instr_rdata_c_id [13]),
    .A1(net650),
    .S(net834),
    .X(\i_ibex/if_stage_i/_040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout550 (.A(net551),
    .X(net550),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_784_  (.A0(\i_ibex/instr_rdata_c_id [14]),
    .A1(net662),
    .S(net831),
    .X(\i_ibex/if_stage_i/_041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_785_  (.A0(\i_ibex/instr_rdata_c_id [15]),
    .A1(net669),
    .S(net832),
    .X(\i_ibex/if_stage_i/_042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_786_  (.A0(\i_ibex/instr_rdata_c_id [1]),
    .A1(net1343),
    .S(net829),
    .X(\i_ibex/if_stage_i/_043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_787_  (.A0(\i_ibex/instr_rdata_c_id [2]),
    .A1(net1350),
    .S(net830),
    .X(\i_ibex/if_stage_i/_044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_788_  (.A0(\i_ibex/instr_rdata_c_id [3]),
    .A1(net1351),
    .S(net829),
    .X(\i_ibex/if_stage_i/_045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_789_  (.A0(\i_ibex/instr_rdata_c_id [4]),
    .A1(net1353),
    .S(net830),
    .X(\i_ibex/if_stage_i/_046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_790_  (.A0(\i_ibex/instr_rdata_c_id [5]),
    .A1(net641),
    .S(net831),
    .X(\i_ibex/if_stage_i/_047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_791_  (.A0(\i_ibex/instr_rdata_c_id [6]),
    .A1(\i_ibex/if_stage_i/fetch_rdata [6]),
    .S(net831),
    .X(\i_ibex/if_stage_i/_048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_792_  (.A0(\i_ibex/instr_rdata_c_id [7]),
    .A1(net1354),
    .S(net830),
    .X(\i_ibex/if_stage_i/_049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_793_  (.A0(\i_ibex/instr_rdata_c_id [8]),
    .A1(net642),
    .S(net830),
    .X(\i_ibex/if_stage_i/_050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout549 (.A(\i_ibex/alu_operand_a_ex [6]),
    .X(net549),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_795_  (.A0(\i_ibex/instr_rdata_c_id [9]),
    .A1(net1357),
    .S(net830),
    .X(\i_ibex/if_stage_i/_051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/_796_  (.Y(\i_ibex/if_stage_i/_352_ ),
    .B(\i_ibex/instr_valid_id ),
    .A_N(\i_ibex/instr_valid_clear ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/_797_  (.B1(\i_ibex/if_stage_i/_352_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_valid_id_d ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/_339_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_798_  (.A0(\i_ibex/pc_id [0]),
    .A1(net380),
    .S(net837),
    .X(\i_ibex/if_stage_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_799_  (.A0(\i_ibex/pc_id [10]),
    .A1(\i_ibex/pc_if [10]),
    .S(net837),
    .X(\i_ibex/if_stage_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_800_  (.A0(\i_ibex/pc_id [11]),
    .A1(\i_ibex/pc_if [11]),
    .S(net837),
    .X(\i_ibex/if_stage_i/_054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_801_  (.A0(\i_ibex/pc_id [12]),
    .A1(\i_ibex/pc_if [12]),
    .S(net837),
    .X(\i_ibex/if_stage_i/_055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_802_  (.A0(\i_ibex/pc_id [13]),
    .A1(\i_ibex/pc_if [13]),
    .S(net842),
    .X(\i_ibex/if_stage_i/_056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_803_  (.A0(\i_ibex/pc_id [14]),
    .A1(\i_ibex/pc_if [14]),
    .S(net842),
    .X(\i_ibex/if_stage_i/_057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_804_  (.A0(\i_ibex/pc_id [15]),
    .A1(\i_ibex/pc_if [15]),
    .S(net842),
    .X(\i_ibex/if_stage_i/_058_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_805_  (.A0(\i_ibex/pc_id [16]),
    .A1(\i_ibex/pc_if [16]),
    .S(net844),
    .X(\i_ibex/if_stage_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_806_  (.A0(\i_ibex/pc_id [17]),
    .A1(\i_ibex/pc_if [17]),
    .S(net844),
    .X(\i_ibex/if_stage_i/_060_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_808_  (.A0(\i_ibex/pc_id [18]),
    .A1(\i_ibex/pc_if [18]),
    .S(net844),
    .X(\i_ibex/if_stage_i/_061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_809_  (.A0(\i_ibex/pc_id [19]),
    .A1(\i_ibex/pc_if [19]),
    .S(net844),
    .X(\i_ibex/if_stage_i/_062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_810_  (.A0(\i_ibex/pc_id [1]),
    .A1(net1478),
    .S(net841),
    .X(\i_ibex/if_stage_i/_063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_811_  (.A0(\i_ibex/pc_id [20]),
    .A1(\i_ibex/pc_if [20]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_064_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_812_  (.A0(\i_ibex/pc_id [21]),
    .A1(\i_ibex/pc_if [21]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_813_  (.A0(\i_ibex/pc_id [22]),
    .A1(\i_ibex/pc_if [22]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_066_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_814_  (.A0(\i_ibex/pc_id [23]),
    .A1(\i_ibex/pc_if [23]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_067_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_815_  (.A0(\i_ibex/pc_id [24]),
    .A1(\i_ibex/pc_if [24]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_816_  (.A0(\i_ibex/pc_id [25]),
    .A1(\i_ibex/pc_if [25]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_817_  (.A0(\i_ibex/pc_id [26]),
    .A1(\i_ibex/pc_if [26]),
    .S(net843),
    .X(\i_ibex/if_stage_i/_070_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout547 (.A(\i_ibex/alu_operand_a_ex [5]),
    .X(net547),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_819_  (.A0(\i_ibex/pc_id [27]),
    .A1(\i_ibex/pc_if [27]),
    .S(net842),
    .X(\i_ibex/if_stage_i/_071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_820_  (.A0(\i_ibex/pc_id [28]),
    .A1(\i_ibex/pc_if [28]),
    .S(net845),
    .X(\i_ibex/if_stage_i/_072_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_821_  (.A0(\i_ibex/pc_id [29]),
    .A1(\i_ibex/pc_if [29]),
    .S(net842),
    .X(\i_ibex/if_stage_i/_073_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_822_  (.A0(\i_ibex/pc_id [2]),
    .A1(\i_ibex/pc_if [2]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_823_  (.A0(\i_ibex/pc_id [30]),
    .A1(\i_ibex/pc_if [30]),
    .S(net844),
    .X(\i_ibex/if_stage_i/_075_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_824_  (.A0(\i_ibex/pc_id [31]),
    .A1(\i_ibex/pc_if [31]),
    .S(net845),
    .X(\i_ibex/if_stage_i/_076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_825_  (.A0(\i_ibex/pc_id [3]),
    .A1(\i_ibex/pc_if [3]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_826_  (.A0(\i_ibex/pc_id [4]),
    .A1(\i_ibex/pc_if [4]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_827_  (.A0(\i_ibex/pc_id [5]),
    .A1(\i_ibex/pc_if [5]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_828_  (.A0(\i_ibex/pc_id [6]),
    .A1(\i_ibex/pc_if [6]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_829_  (.A0(\i_ibex/pc_id [7]),
    .A1(\i_ibex/pc_if [7]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_830_  (.A0(\i_ibex/pc_id [8]),
    .A1(\i_ibex/pc_if [8]),
    .S(net842),
    .X(\i_ibex/if_stage_i/_082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/_831_  (.A0(\i_ibex/pc_id [9]),
    .A1(\i_ibex/pc_if [9]),
    .S(net841),
    .X(\i_ibex/if_stage_i/_083_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/cs_registers_i/_2511__379  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net379));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_440_  (.A(net644),
    .B(net1358),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_407_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout545 (.A(\i_ibex/alu_operand_a_ex [4]),
    .X(net545),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_443_  (.A(net1357),
    .B(net643),
    .C(net1354),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_410_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_444_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_411_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_407_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_410_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout543 (.A(\i_ibex/alu_operand_a_ex [3]),
    .X(net543),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_447_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_414_ ),
    .A(net669),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_448_  (.A(net647),
    .B(net1326),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_415_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout541 (.A(\i_ibex/alu_operand_a_ex [2]),
    .X(net541),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout539 (.A(\i_ibex/alu_operand_a_ex [28]),
    .X(net539),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_453_  (.A(net641),
    .B(\i_ibex/if_stage_i/fetch_rdata [6]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_420_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout538 (.A(net539),
    .X(net538),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout537 (.A(\i_ibex/alu_operand_a_ex [1]),
    .X(net537),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_456_  (.A(net1353),
    .B(net1351),
    .C(net1350),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_423_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_457_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_424_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_420_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_423_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_459_  (.A(net659),
    .B(net1274),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_426_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/if_stage_i/compressed_decoder_i/_460_  (.A(net671),
    .B_N(net658),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_427_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_461_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_415_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_426_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_428_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_427_ ));
 sg13g2_buf_2 fanout535 (.A(\i_ibex/alu_operand_a_ex [0]),
    .X(net535),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout534 (.A(\i_ibex/alu_operand_a_ex [27]),
    .X(net534),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_464_  (.A(net667),
    .B(net662),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_431_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_466_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_433_ ),
    .A(net650),
    .VSS(VSS));
 sg13g2_buf_2 fanout532 (.A(\i_ibex/alu_operand_a_ex [26]),
    .X(net532),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout531 (.A(net532),
    .X(net531),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_469_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_436_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_433_ ),
    .B(net1347),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_470_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net649),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_431_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_437_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_436_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_471_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_437_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_438_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_411_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_428_ ));
 sg13g2_buf_2 fanout530 (.A(\i_ibex/alu_operand_a_ex [25]),
    .X(net530),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/if_stage_i/compressed_decoder_i/_473_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_000_ ),
    .B(net650),
    .A(net669));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/if_stage_i/compressed_decoder_i/_475_  (.A(net647),
    .B(net641),
    .C(\i_ibex/if_stage_i/fetch_rdata [6]),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_411_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_476_  (.A(net1347),
    .B(net1284),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_002_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_477_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_004_ ),
    .A(net663),
    .B(net1287),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_478_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_005_ ),
    .A(net636),
    .VSS(VSS));
 sg13g2_buf_2 fanout528 (.A(\i_ibex/alu_operand_a_ex [24]),
    .X(net528),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_480_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_005_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_007_ ),
    .VSS(VSS),
    .A1(net1347),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_004_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_481_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_003_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_007_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/if_stage_i/compressed_decoder_i/_483_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .A(net1358),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_484_  (.A(net662),
    .B_N(net667),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_485_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ),
    .A(net1287),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_486_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net645),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_013_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ));
 sg13g2_buf_2 fanout526 (.A(\i_ibex/alu_operand_b_ex [1]),
    .X(net526),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 load_slew525 (.A(net1140),
    .X(net525),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_489_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_016_ ),
    .A(net654),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_427_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_490_  (.A(net647),
    .B(net1274),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_016_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_491_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net649),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_013_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_018_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_017_ ));
 sg13g2_nand2b_2 \i_ibex/if_stage_i/compressed_decoder_i/_492_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_019_ ),
    .B(net638),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1343));
 sg13g2_buf_1 max_cap524 (.A(net1130),
    .X(net524),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_494_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_018_ ),
    .B(net1323),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_495_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_008_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_438_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_021_ ),
    .X(\i_ibex/if_stage_i/illegal_c_insn ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/if_stage_i/compressed_decoder_i/_496_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ),
    .B(net669),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net658));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_497_  (.B1(net1285),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_023_ ),
    .VSS(VSS),
    .A1(net1343),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_498_  (.Y(\i_ibex/if_stage_i/instr_decompressed [0]),
    .A(net626),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_499_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_024_ ),
    .A(net1343),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_500_  (.A(net1322),
    .B(net626),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 \i_ibex/if_stage_i/compressed_decoder_i/_501_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_025_ ),
    .Y(\i_ibex/if_stage_i/instr_is_compressed ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_502_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .A(\i_ibex/if_stage_i/instr_decompressed [0]),
    .B(\i_ibex/if_stage_i/instr_is_compressed ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_503_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_027_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [31]),
    .B(net644),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_504_  (.A(net1345),
    .B(net626),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 load_slew523 (.A(net1125),
    .X(net523),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_506_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_030_ ),
    .A(net649),
    .B(net1282),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_507_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_013_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_027_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_031_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_030_ ));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_508_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [31]),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_031_ ),
    .X(\i_ibex/if_stage_i/instr_decompressed [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_509_  (.B(net645),
    .C(net1358),
    .A(net648),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(\i_ibex/csr_addr [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_511_  (.A(\i_ibex/if_stage_i/fetch_rdata [30]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_032_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net522),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net521),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_514_  (.B1(net670),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_037_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_407_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_034_ ));
 sg13g2_inv_2 \i_ibex/if_stage_i/compressed_decoder_i/_515_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .A(net646),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_516_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_039_ ),
    .A(net644),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_517_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_518_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_040_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_041_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_039_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_420_ ));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net521),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout518 (.A(net521),
    .X(net518),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_521_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_041_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_044_ ),
    .B1(net652));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_522_  (.A(net658),
    .B(net1286),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout517 (.A(net522),
    .X(net517),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_524_  (.A(net646),
    .B(net663),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_525_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net642),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_047_ ),
    .B1(net1273),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_037_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_048_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_044_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_526_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_049_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [30]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_527_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_049_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [30]),
    .VSS(VSS),
    .A1(net1323),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_048_ ));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_528_  (.A(net658),
    .B(net654),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_529_  (.A(net1357),
    .B(net1355),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_530_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_407_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_051_ ),
    .A(net642),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/if_stage_i/compressed_decoder_i/_531_  (.A(net646),
    .B(net658),
    .C(net650),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout516 (.A(net522),
    .X(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_533_  (.B1(net1325),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_055_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_053_ ));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(net522),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_536_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net669),
    .A2(net1280),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_058_ ),
    .B1(net651));
 sg13g2_nor2b_2 \i_ibex/if_stage_i/compressed_decoder_i/_537_  (.A(net654),
    .B_N(net659),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_538_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_060_ ),
    .A(net1325),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_539_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_060_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_061_ ),
    .VSS(VSS),
    .A1(net661),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_058_ ));
 sg13g2_nor4_2 \i_ibex/if_stage_i/compressed_decoder_i/_540_  (.A(net1325),
    .B(net659),
    .C(net654),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_062_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net1280));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_541_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_063_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_062_ ),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_542_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_064_ ),
    .A(net1322),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_543_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/fetch_rdata [21]),
    .C1(net625),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_064_ ),
    .A1(net1351),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_065_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_061_ ));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(net515),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(net515),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_546_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_068_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [21]),
    .VSS(VSS));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(net515),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_548_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_070_ ),
    .A(net1285),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_431_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_549_  (.A(net1351),
    .B(net1345),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_070_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_550_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_068_ ),
    .A2(net1345),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_072_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_071_ ));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net515),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_552_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_074_ ),
    .A(net672),
    .B(net658),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_553_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_074_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_075_ ),
    .VSS(VSS),
    .A1(net659),
    .A2(net1322));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net515),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_555_  (.A(net656),
    .B_N(net1351),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_556_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_078_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_075_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_077_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_023_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_557_  (.A(net637),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_078_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_558_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net639),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_072_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_080_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_079_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_559_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_055_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_065_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [21]),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_080_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_560_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1285),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_081_ ),
    .B1(net1344));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_561_  (.A(net625),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_081_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_562_  (.B1(\i_ibex/if_stage_i/fetch_rdata [20]),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_083_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_025_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_082_ ));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_563_  (.A(net1345),
    .B(net638),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/compressed_decoder_i/_565_  (.B(net1350),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .A(net671),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_086_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(net620));
 sg13g2_and3_1 \i_ibex/if_stage_i/compressed_decoder_i/_566_  (.X(\i_ibex/if_stage_i/compressed_decoder_i/_087_ ),
    .A(net646),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_407_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_410_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_567_  (.A(net1274),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_568_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_089_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [2]),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_569_  (.A(net653),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_089_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_427_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_090_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_570_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_088_ ),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_090_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_087_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [20]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_091_ ),
    .A2(net655));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_571_  (.A(net1322),
    .B(net638),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_572_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_093_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .A_N(\i_ibex/if_stage_i/compressed_decoder_i/_091_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/if_stage_i/compressed_decoder_i/_573_  (.X(\i_ibex/if_stage_i/compressed_decoder_i/_094_ ),
    .A(net642),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_407_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_574_  (.B1(net663),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_095_ ),
    .VSS(VSS),
    .A1(net672),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_094_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_575_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [12]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_095_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_096_ ),
    .B1(net1286));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_576_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_097_ ),
    .A(net1350),
    .B(net1280),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/if_stage_i/compressed_decoder_i/_577_  (.X(\i_ibex/if_stage_i/compressed_decoder_i/_098_ ),
    .A(net646),
    .B(net644),
    .C(net1359),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_578_  (.B(net669),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_098_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [20]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_099_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_579_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_097_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_099_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_100_ ),
    .B1(net659));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_580_  (.A(net668),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_089_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_581_  (.A(net652),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_100_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_101_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/if_stage_i/compressed_decoder_i/_582_  (.A(net1324),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_096_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_102_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/compressed_decoder_i/_583_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_086_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_093_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_083_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [20]),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_103_ ));
 sg13g2_nor3_2 \i_ibex/if_stage_i/compressed_decoder_i/_584_  (.A(net667),
    .B(net662),
    .C(net654),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_585_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_105_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_039_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_586_  (.A(net651),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_011_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_587_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_107_ ),
    .A(net1322),
    .B(net625),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_588_  (.B1(\i_ibex/if_stage_i/instr_is_compressed ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_108_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_106_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_107_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_589_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_109_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_108_ ),
    .B2(\i_ibex/if_stage_i/fetch_rdata [19]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_105_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_590_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_110_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .B(net1275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_591_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_039_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_593_  (.A(net667),
    .B(net654),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_594_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [19]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_084_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_114_ ),
    .B1(net1272));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_595_  (.B1(\i_ibex/if_stage_i/fetch_rdata [19]),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_115_ ),
    .VSS(VSS),
    .A1(net652),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_025_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_596_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_115_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_116_ ),
    .VSS(VSS),
    .A1(net661),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_114_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_597_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_110_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_111_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_117_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_116_ ));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_599_  (.A(net644),
    .B(net1359),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_600_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [19]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_119_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_120_ ),
    .B1(net651));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_601_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_121_ ),
    .B(\i_ibex/if_stage_i/fetch_rdata [12]),
    .A_N(\i_ibex/if_stage_i/compressed_decoder_i/_120_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_602_  (.B(net652),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ),
    .A(net1326),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_603_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_123_ ),
    .A(net1281),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_604_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net661),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_123_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_122_ ),
    .A1(net1283),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_124_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_121_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_605_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_125_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_124_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_606_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_125_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [19]),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_109_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_117_ ));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_607_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_126_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [12]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_608_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_127_ ),
    .B(net1359),
    .A_N(net658),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_609_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1272),
    .C1(net1324),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_127_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_128_ ),
    .A2(net1273));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_610_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_128_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_129_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/fetch_rdata [18]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_063_ ));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_611_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_126_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_427_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_129_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_612_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_131_ ),
    .A(net1285),
    .B(net625),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_613_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_131_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [18]),
    .B1(net1322),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_132_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_614_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_133_ ),
    .B(net669),
    .A_N(net646),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_615_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_133_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_423_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_134_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_616_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_135_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_133_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_420_ ));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_617_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_134_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_135_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_618_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_137_ ),
    .A(net1345),
    .B(net625),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_619_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_137_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_138_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_620_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_139_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_136_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_138_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_132_ ),
    .A1(net1324),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_621_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/fetch_rdata [18]),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_107_ ),
    .B1(net1283),
    .A1(net664),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_140_ ),
    .A2(net1285));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_622_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_130_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_139_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [18]),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_140_ ));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_624_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_142_ ),
    .B1(net1356),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_136_ ),
    .A2(net656),
    .A1(\i_ibex/if_stage_i/fetch_rdata [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_625_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_143_ ),
    .A(net648),
    .B(net650),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_626_  (.B(net663),
    .C(net1356),
    .A(net672),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_627_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_144_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_145_ ),
    .VSS(VSS),
    .A1(net659),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_143_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_628_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_146_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [17]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_629_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_147_ ),
    .A(net1356),
    .B(net1280),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_630_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_146_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_147_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_148_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_631_  (.A(\i_ibex/if_stage_i/fetch_rdata [17]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_025_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_149_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/if_stage_i/compressed_decoder_i/_632_  (.A(net620),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_145_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_148_ ),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_149_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_633_  (.B1(net638),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_151_ ),
    .VSS(VSS),
    .A1(net1356),
    .A2(net1283));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_634_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_152_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_151_ ),
    .A_N(net659),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_635_  (.A(net655),
    .B_N(net1356),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_153_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_636_  (.A(net637),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_153_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_637_  (.A(net1345),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_154_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_638_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_156_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_152_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_155_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_108_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_639_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_150_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_055_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_156_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_640_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_157_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [17]),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_137_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_142_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_641_  (.A(net642),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_098_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_642_  (.A(net652),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_643_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_159_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_160_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/fetch_rdata [16]),
    .A2(net1280));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_644_  (.A(net668),
    .B(net662),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/if_stage_i/compressed_decoder_i/_645_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_646_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_163_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 \i_ibex/if_stage_i/compressed_decoder_i/_647_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_164_ ),
    .B(net662),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net667));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_648_  (.A(net1287),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_164_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_650_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1284),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_143_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_167_ ),
    .B1(net665));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_651_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_165_ ),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_167_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_163_ ),
    .A1(net643),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_168_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_161_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_652_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_168_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_169_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_158_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_160_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_653_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_170_ ),
    .A(net642),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_654_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_170_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_104_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_171_ ),
    .B1(net1324));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_655_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_172_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [16]),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_656_  (.A(net650),
    .B(net643),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_173_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_657_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_172_ ),
    .A2(net654),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_174_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_173_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_658_  (.B(net1274),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_415_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_659_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_176_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_174_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_175_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_660_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [16]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_025_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_177_ ),
    .B1(net620));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_661_  (.A(\i_ibex/if_stage_i/fetch_rdata [16]),
    .B(net636),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_662_  (.B1(net1324),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_179_ ),
    .VSS(VSS),
    .A1(net1322),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_178_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_663_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_180_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_179_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_431_ ),
    .A2(net620),
    .A1(net662),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_664_  (.B(net1283),
    .C(net620),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_172_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_181_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_665_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_181_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_182_ ),
    .VSS(VSS),
    .A1(net652),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_180_ ));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_667_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_172_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_184_ ),
    .VSS(VSS),
    .A1(net636),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_081_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_668_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_185_ ),
    .A(net1324),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_669_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_170_ ),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_185_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_182_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_176_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_186_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_177_ ));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_670_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_171_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_169_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_186_ ),
    .X(\i_ibex/if_stage_i/instr_decompressed [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/if_stage_i/compressed_decoder_i/_671_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_016_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_094_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 \i_ibex/if_stage_i/compressed_decoder_i/_673_  (.A(net654),
    .B_N(net667),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_674_  (.A(net1355),
    .B_N(\i_ibex/if_stage_i/compressed_decoder_i/_189_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_675_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_191_ ),
    .A(net671),
    .B(net1355),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_676_  (.A(net647),
    .B(net666),
    .C(net1287),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_677_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net661),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_192_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_191_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_032_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_193_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_190_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_678_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [5]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_187_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_194_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_193_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_679_  (.B1(net1281),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_195_ ),
    .VSS(VSS),
    .A1(net1354),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_070_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_680_  (.A(net1325),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_681_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1354),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_197_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_196_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_682_  (.A(net650),
    .B(net638),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_683_  (.B1(net1345),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_199_ ),
    .VSS(VSS),
    .A1(net1325),
    .A2(net1279));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_684_  (.A(net639),
    .B_N(net1354),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_685_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_201_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_200_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_136_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_199_ ),
    .A1(net1324),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_686_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_197_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_084_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_201_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_687_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_202_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [15]),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_194_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_195_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_688_  (.A(net1323),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_104_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_689_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_187_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_203_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [4]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_690_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_019_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_131_ ),
    .A(net664),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_691_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_119_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_206_ ),
    .VSS(VSS),
    .A1(net647),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_420_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_692_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_207_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_189_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_206_ ),
    .A2(net656),
    .A1(net647),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 \i_ibex/if_stage_i/compressed_decoder_i/_693_  (.A(net664),
    .B(net1323),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_207_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_208_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_694_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_205_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_208_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_204_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_695_  (.B1(net1359),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_209_ ),
    .VSS(VSS),
    .A1(net647),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_696_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_209_ ),
    .C1(net1323),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_111_ ),
    .A1(net649),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_210_ ),
    .A2(net1273));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_697_  (.A2(net639),
    .A1(net671),
    .B1(net663),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_698_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/instr_is_compressed ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_211_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_212_ ),
    .B1(net653));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_699_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_213_ ),
    .A(net1352),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_187_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_700_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_213_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [13]),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_210_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_212_ ));
 sg13g2_nand2_2 \i_ibex/if_stage_i/compressed_decoder_i/_701_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .A(net1285),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_702_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net649),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_215_ ),
    .B1(net636));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_703_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_216_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_104_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_704_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_216_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_217_ ),
    .VSS(VSS),
    .A1(net1349),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_215_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_705_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_218_ ),
    .A(net645),
    .B(net1358),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_706_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [5]),
    .A2(\i_ibex/if_stage_i/fetch_rdata [6]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_219_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_218_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_707_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_220_ ),
    .VSS(VSS),
    .A1(net651),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_219_ ));
 sg13g2_nand3b_1 \i_ibex/if_stage_i/compressed_decoder_i/_708_  (.B(net1284),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_220_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_221_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net665));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_709_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_222_ ),
    .A(net656),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_710_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_221_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_222_ ),
    .A(net639),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_711_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_224_ ),
    .A(net648),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_712_  (.B(net1281),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_187_ ),
    .A(net1350),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_714_  (.A(net1322),
    .B(net1279),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_715_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_228_ ),
    .A(net648),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_716_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_229_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_225_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_228_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_224_ ),
    .A1(net620),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_717_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_223_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_217_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_229_ ),
    .X(\i_ibex/if_stage_i/instr_decompressed [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(net517),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_719_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_231_ ),
    .A(net648),
    .B(net637),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_720_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_231_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_232_ ),
    .VSS(VSS),
    .A1(net636),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_127_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_721_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_233_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_232_ ),
    .B2(net1272),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_047_ ),
    .A1(net637),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/compressed_decoder_i/_722_  (.B(net670),
    .C(net644),
    .A(net648),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_723_  (.A(\i_ibex/if_stage_i/fetch_rdata [29]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_235_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_724_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_236_ ),
    .A(net1358),
    .B(net1273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_725_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_236_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_237_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_235_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_726_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_238_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_203_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_237_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_727_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_238_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [29]),
    .VSS(VSS),
    .A1(net1347),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_233_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_728_  (.A(net668),
    .B(net1348),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_239_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/if_stage_i/compressed_decoder_i/_729_  (.A(net1326),
    .B(net666),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_024_ ),
    .D(net1275),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_240_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_730_  (.B1(net1278),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_241_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_239_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_240_ ));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_731_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_242_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_203_ ),
    .A_N(net661),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_732_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_241_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_242_ ),
    .A(net645),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_243_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_733_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_243_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [11]),
    .VSS(VSS),
    .A1(net1324),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_063_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_734_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_244_ ),
    .VSS(VSS),
    .A1(net625),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_022_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_735_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .A2(net1283),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_245_ ),
    .B1(net636));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_736_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1285),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_245_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_244_ ),
    .A1(net664),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_246_ ),
    .A2(net1359));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_737_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_247_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_005_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_738_  (.B(net1344),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_247_ ),
    .A(net1359),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_248_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_739_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_248_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [10]),
    .VSS(VSS),
    .A1(net1343),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_246_ ));
 sg13g2_inv_2 \i_ibex/if_stage_i/compressed_decoder_i/_740_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_249_ ),
    .A(net1353),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_741_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_250_ ),
    .A(net1356),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/compressed_decoder_i/_742_  (.A0(\i_ibex/if_stage_i/compressed_decoder_i/_249_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_250_ ),
    .S(net1325),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_743_  (.A(net661),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_153_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_252_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_744_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net664),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_251_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_253_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_252_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_745_  (.B(net670),
    .C(net660),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_746_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_254_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_255_ ),
    .VSS(VSS),
    .A1(net668),
    .A2(net1353));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_747_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1285),
    .C1(net636),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_255_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_250_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_256_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_748_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net639),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_253_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_257_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_256_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_749_  (.B(net1356),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_247_ ),
    .A(net1343),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_750_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_258_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [9]),
    .VSS(VSS),
    .A1(net1343),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_257_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_751_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_259_ ),
    .A(net1286),
    .B(net642),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_752_  (.B(net1351),
    .C(net637),
    .A(net663),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_753_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_260_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_261_ ),
    .VSS(VSS),
    .A1(net660),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_259_ ));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_754_  (.A(net639),
    .B_N(net1351),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_755_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_263_ ),
    .B(net651),
    .A_N(net660),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_756_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1325),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_263_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_264_ ),
    .B1(net625));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_757_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_170_ ),
    .B(net1279),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_264_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_265_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_758_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1272),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_265_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_262_ ),
    .A1(net671),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_266_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_261_ ));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_759_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_267_ ),
    .B(net1275),
    .A_N(net665),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_760_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_189_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_267_ ),
    .A(net626),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_761_  (.B(net643),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_268_ ),
    .A(net1346),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_269_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_762_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_269_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [8]),
    .VSS(VSS),
    .A1(net1346),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_266_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_763_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_270_ ),
    .A(net649),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_411_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_764_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_271_ ),
    .A(net1355),
    .B(net1274),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_765_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_271_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_272_ ),
    .VSS(VSS),
    .A1(net1274),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_270_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_766_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_272_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_159_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_273_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_767_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_189_ ),
    .B_N(net1354),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_274_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_768_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_275_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .B(net660),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_769_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_276_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_263_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_275_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_770_  (.B(net1281),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_276_ ),
    .A(net671),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_277_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_771_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_278_ ),
    .A(net638),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_772_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1325),
    .A2(net1273),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_279_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_278_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_773_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_280_ ),
    .A(net639),
    .B(net1354),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_774_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_280_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_281_ ),
    .VSS(VSS),
    .A1(net1345),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_279_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_775_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_282_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_277_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_281_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_274_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_776_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1354),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_107_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .A1(net1350),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_283_ ),
    .A2(net1272));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_777_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_273_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_282_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [7]),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_283_ ));
 sg13g2_nor4_1 \i_ibex/if_stage_i/compressed_decoder_i/_778_  (.A(net660),
    .B(net651),
    .C(net1275),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_137_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_284_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_779_  (.A(net658),
    .B(net1281),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_285_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_780_  (.B1(net670),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_286_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_284_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_285_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_781_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_287_ ),
    .A(net1282),
    .B(net1273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_782_  (.A(net1348),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ),
    .C(net1280),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_288_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_783_  (.B1(\i_ibex/if_stage_i/fetch_rdata [6]),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_289_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_288_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_784_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_287_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_289_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_286_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_785_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_290_ ),
    .A(net641),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_786_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net648),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_290_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_291_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_218_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_787_  (.B1(net669),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_292_ ),
    .VSS(VSS),
    .A1(net661),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_291_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_788_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_293_ ),
    .A(net1287),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_292_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_789_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_293_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_294_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_164_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_790_  (.A(net661),
    .B(net1348),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_791_  (.B1(net626),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_296_ ),
    .VSS(VSS),
    .A1(net653),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_295_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_792_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/instr_is_compressed ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_296_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_297_ ),
    .B1(net641));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_793_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1282),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_297_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_294_ ),
    .A1(net1326),
    .Y(\i_ibex/if_stage_i/instr_decompressed [5]),
    .A2(net1278));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_794_  (.B1(net1347),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_298_ ),
    .VSS(VSS),
    .A1(net1274),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_087_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_795_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_299_ ),
    .A(net626),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_796_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net670),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_298_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_300_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_299_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_797_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net670),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_098_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_301_ ),
    .B1(net1347));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_798_  (.B1(net626),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_302_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_249_ ),
    .A2(net1343));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_799_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_303_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_800_  (.B1(net639),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_304_ ),
    .VSS(VSS),
    .A1(net1344),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_427_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_801_  (.B(net1353),
    .C(net625),
    .A(net655),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_802_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_304_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_305_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_303_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_306_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_803_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_306_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_307_ ),
    .VSS(VSS),
    .A1(net1353),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_301_ ));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_804_  (.Y(\i_ibex/if_stage_i/instr_decompressed [4]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_307_ ),
    .A_N(\i_ibex/if_stage_i/compressed_decoder_i/_300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_805_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1352),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_062_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_308_ ),
    .B1(net1273));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_806_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_309_ ),
    .A(net1352),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_807_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_309_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [3]),
    .VSS(VSS),
    .A1(net1323),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_308_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_808_  (.B1(net638),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_310_ ),
    .VSS(VSS),
    .A1(net651),
    .A2(net1280));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_809_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_310_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_311_ ),
    .B1(net1344));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_810_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_089_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_092_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_311_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_811_  (.A(net1274),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_012_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_087_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_812_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net655),
    .A2(net1350),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_314_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_313_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_813_  (.B(net1281),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_095_ ),
    .A(net656),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_814_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_315_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_316_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_137_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_314_ ));
 sg13g2_or2_1 \i_ibex/if_stage_i/compressed_decoder_i/_815_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/instr_decompressed [2]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_316_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_312_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_816_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_126_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_317_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_249_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_817_  (.B(net1282),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_317_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_165_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_318_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_818_  (.A(net646),
    .B(net671),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/compressed_decoder_i/_819_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1323),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_320_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_319_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_820_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_321_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_320_ ),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_821_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_321_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_822_  (.B1(\i_ibex/if_stage_i/fetch_rdata [28]),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_323_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_026_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_322_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_823_  (.A(net1358),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_324_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_824_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net655),
    .A2(net1357),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_325_ ),
    .B1(net1272));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_825_  (.B1(net649),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_326_ ),
    .VSS(VSS),
    .A1(net1272),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_161_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_826_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_326_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_327_ ),
    .VSS(VSS),
    .A1(net660),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_325_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_827_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_320_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_328_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_324_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_327_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_828_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_104_ ),
    .C(net620),
    .A(net1356),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/compressed_decoder_i/_829_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_323_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_328_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_318_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [28]),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_329_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_830_  (.Y(\i_ibex/if_stage_i/instr_decompressed [1]),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_081_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_831_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_016_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_094_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_832_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net649),
    .A2(net1287),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_331_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_164_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_833_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net668),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_331_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_050_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_332_ ),
    .A2(net1284));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_834_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .B(\i_ibex/if_stage_i/fetch_rdata [27]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_333_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_835_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_165_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_094_ ),
    .A(net1352),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_334_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_836_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_334_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_335_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_333_ ));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_837_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_330_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_332_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_335_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_838_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_170_ ),
    .B(net1283),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_337_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_839_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [27]),
    .A2(net1284),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_338_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_337_ ));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_840_  (.A(net637),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_338_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_339_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_841_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_340_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [27]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/compressed_decoder_i/_842_  (.A0(net1351),
    .A1(net642),
    .S(net667),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_341_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_843_  (.B(net1278),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_341_ ),
    .A(net663),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_342_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_844_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_340_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_342_ ),
    .A(net1348),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_845_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_343_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_344_ ),
    .VSS(VSS),
    .A1(net1348),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_339_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_846_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_344_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/instr_decompressed [27]),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_321_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_336_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_847_  (.B1(net1326),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_345_ ),
    .VSS(VSS),
    .A1(net1287),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_848_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_285_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_345_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [5]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_346_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_849_  (.A(net668),
    .B(net666),
    .C(net1355),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_347_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_850_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_290_ ),
    .A2(net664),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_348_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_347_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_851_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_084_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_349_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/fetch_rdata [26]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_106_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_852_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_350_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_349_ ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_853_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_350_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_351_ ),
    .VSS(VSS),
    .A1(net653),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_348_ ));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_854_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_101_ ),
    .B_N(\i_ibex/if_stage_i/compressed_decoder_i/_191_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_352_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_855_  (.A(net637),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_004_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_352_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_353_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/compressed_decoder_i/_856_  (.A(net1278),
    .B_N(\i_ibex/if_stage_i/fetch_rdata [26]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_354_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_857_  (.B1(net1348),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_355_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_353_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_354_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_858_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_010_ ),
    .B(\i_ibex/if_stage_i/fetch_rdata [26]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_356_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_859_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_357_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_275_ ),
    .B2(net1272),
    .A2(net1273),
    .A1(net1355),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_860_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_357_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_358_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_356_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_861_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_320_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_359_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_330_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_358_ ));
 sg13g2_nand4_1 \i_ibex/if_stage_i/compressed_decoder_i/_862_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_351_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_355_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_346_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [26]),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/compressed_decoder_i/_359_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_863_  (.B1(net1350),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_360_ ),
    .VSS(VSS),
    .A1(net659),
    .A2(net652));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_864_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net668),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_331_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_360_ ),
    .A1(net655),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_361_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_089_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_865_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_362_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [25]),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_866_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1358),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_362_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_363_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_234_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_867_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_320_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_364_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_361_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_363_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_868_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_365_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_047_ ),
    .B(net1278),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_869_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_365_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_366_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_362_ ),
    .A2(net1278));
 sg13g2_mux2_1 \i_ibex/if_stage_i/compressed_decoder_i/_870_  (.A0(\i_ibex/if_stage_i/compressed_decoder_i/_038_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_362_ ),
    .S(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_367_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_871_  (.A(net1347),
    .B(net638),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_367_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_368_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_872_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1347),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_366_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_369_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_368_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_873_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_126_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_370_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_089_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_052_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_874_  (.B(net1282),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_370_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_165_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_371_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_875_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_369_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_371_ ),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_364_ ),
    .Y(\i_ibex/if_stage_i/instr_decompressed [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_876_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_131_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_877_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [24]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_131_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_373_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_372_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_878_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_374_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [6]),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_094_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_879_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_374_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_126_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_016_ ),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_375_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_880_  (.B1(net670),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_376_ ),
    .VSS(VSS),
    .A1(net660),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_119_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_881_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .B(net655),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_377_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_882_  (.B1(net1281),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_378_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_039_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_263_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_883_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_377_ ),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_378_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_376_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [24]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_379_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_062_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_884_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/fetch_rdata [24]),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_107_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_214_ ),
    .A1(net644),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_380_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_113_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_885_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_379_ ),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_380_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_375_ ),
    .A1(net1349),
    .Y(\i_ibex/if_stage_i/instr_decompressed [24]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_373_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/compressed_decoder_i/_886_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_381_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [23]),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_887_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_381_ ),
    .B(net1278),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_382_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_888_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net641),
    .A2(net1278),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_383_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_382_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_889_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net648),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_381_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_384_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_218_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_890_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_385_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_384_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_011_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_376_ ),
    .A1(net641),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/if_stage_i/compressed_decoder_i/_891_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_386_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_385_ ),
    .A(net653));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_892_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net647),
    .C1(net1323),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_187_ ),
    .A1(net641),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_387_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_045_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_893_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_059_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_388_ ),
    .VSS(VSS),
    .A1(net667),
    .A2(net1358));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_894_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_290_ ),
    .B(net662),
    .C(net1283),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_389_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_895_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_rdata [23]),
    .A2(net1283),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_390_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_389_ ));
 sg13g2_and3_1 \i_ibex/if_stage_i/compressed_decoder_i/_896_  (.X(\i_ibex/if_stage_i/compressed_decoder_i/_391_ ),
    .A(net620),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_388_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_897_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_387_ ),
    .C1(\i_ibex/if_stage_i/compressed_decoder_i/_391_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_386_ ),
    .A1(net1349),
    .Y(\i_ibex/if_stage_i/instr_decompressed [23]),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_383_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/compressed_decoder_i/_898_  (.A(net652),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_249_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_392_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/compressed_decoder_i/_899_  (.A0(\i_ibex/if_stage_i/fetch_rdata [22]),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_392_ ),
    .S(net660),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_393_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/compressed_decoder_i/_900_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_394_ ),
    .A(net671),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_393_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/compressed_decoder_i/_901_  (.A(net650),
    .B(\i_ibex/if_stage_i/fetch_rdata [22]),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_395_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_902_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_162_ ),
    .B(net670),
    .C(net656),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_396_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/compressed_decoder_i/_903_  (.A(\i_ibex/if_stage_i/compressed_decoder_i/_107_ ),
    .B(\i_ibex/if_stage_i/compressed_decoder_i/_395_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_396_ ),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_904_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net664),
    .A2(net655),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_398_ ),
    .B1(net1353));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_905_  (.B1(net1353),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_399_ ),
    .VSS(VSS),
    .A1(net651),
    .A2(net1280));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_906_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_098_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_189_ ),
    .A(\i_ibex/if_stage_i/fetch_rdata [22]),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_400_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/compressed_decoder_i/_907_  (.A2(\i_ibex/if_stage_i/compressed_decoder_i/_400_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_399_ ),
    .B1(net664),
    .X(\i_ibex/if_stage_i/compressed_decoder_i/_401_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_908_  (.B1(\i_ibex/if_stage_i/compressed_decoder_i/_401_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_402_ ),
    .VSS(VSS),
    .A1(net668),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_398_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_909_  (.B(net653),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_126_ ),
    .A(net663),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_403_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/compressed_decoder_i/_910_  (.B(\i_ibex/if_stage_i/compressed_decoder_i/_402_ ),
    .C(\i_ibex/if_stage_i/compressed_decoder_i/_403_ ),
    .A(net1281),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_404_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/compressed_decoder_i/_911_  (.B1(net1348),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/compressed_decoder_i/_405_ ),
    .VSS(VSS),
    .A1(net653),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_249_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_912_  (.Y(\i_ibex/if_stage_i/compressed_decoder_i/_406_ ),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_405_ ),
    .B2(net626),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_227_ ),
    .A1(\i_ibex/if_stage_i/fetch_rdata [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/compressed_decoder_i/_913_  (.Y(\i_ibex/if_stage_i/instr_decompressed [22]),
    .B1(\i_ibex/if_stage_i/compressed_decoder_i/_404_ ),
    .B2(\i_ibex/if_stage_i/compressed_decoder_i/_406_ ),
    .A2(\i_ibex/if_stage_i/compressed_decoder_i/_397_ ),
    .A1(\i_ibex/if_stage_i/compressed_decoder_i/_394_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/illegal_c_insn_id_o_reg  (.CLK(clknet_leaf_112_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_000_ ),
    .Q_N(\i_ibex/if_stage_i/_438_ ),
    .Q(\i_ibex/illegal_c_insn_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_fetch_err_o_reg  (.RESET_B(net1577),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_001_ ),
    .Q(\i_ibex/instr_fetch_err ),
    .Q_N(\i_ibex/if_stage_i/_437_ ),
    .CLK(clknet_leaf_89_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_fetch_err_plus2_o_reg  (.RESET_B(net1576),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_002_ ),
    .Q(\i_ibex/instr_fetch_err_plus2 ),
    .Q_N(\i_ibex/if_stage_i/_436_ ),
    .CLK(clknet_leaf_88_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_is_compressed_id_o_reg  (.CLK(clknet_leaf_88_clk_i_regs),
    .RESET_B(net1576),
    .D(\i_ibex/if_stage_i/_003_ ),
    .Q_N(\i_ibex/if_stage_i/_439_ ),
    .Q(\i_ibex/instr_is_compressed_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_new_id_o_reg  (.CLK(clknet_leaf_142_clk_i_regs),
    .RESET_B(net1627),
    .D(net843),
    .Q_N(\i_ibex/if_stage_i/_435_ ),
    .Q(\i_ibex/instr_new_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[0]_reg  (.RESET_B(net1668),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_004_ ),
    .Q(\i_ibex/instr_rdata_id [0]),
    .Q_N(\i_ibex/if_stage_i/_434_ ),
    .CLK(clknet_leaf_112_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[10]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_005_ ),
    .Q(\i_ibex/id_stage_i/imm_s_type [3]),
    .Q_N(\i_ibex/if_stage_i/_433_ ),
    .CLK(clknet_leaf_128_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[11]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_006_ ),
    .Q(\i_ibex/id_stage_i/imm_s_type [4]),
    .Q_N(\i_ibex/if_stage_i/_432_ ),
    .CLK(clknet_leaf_128_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[12]_reg  (.CLK(clknet_leaf_107_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_007_ ),
    .Q_N(\i_ibex/if_stage_i/_431_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[13]_reg  (.CLK(clknet_leaf_111_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_008_ ),
    .Q_N(\i_ibex/if_stage_i/_430_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[14]_reg  (.CLK(clknet_leaf_112_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_009_ ),
    .Q_N(\i_ibex/if_stage_i/_429_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[15]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_010_ ),
    .Q(\i_ibex/id_stage_i/zimm_rs1_type [0]),
    .Q_N(\i_ibex/if_stage_i/_428_ ),
    .CLK(clknet_leaf_129_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[16]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_011_ ),
    .Q(\i_ibex/id_stage_i/zimm_rs1_type [1]),
    .Q_N(\i_ibex/if_stage_i/_427_ ),
    .CLK(clknet_leaf_135_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[17]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_012_ ),
    .Q(\i_ibex/id_stage_i/zimm_rs1_type [2]),
    .Q_N(\i_ibex/if_stage_i/_426_ ),
    .CLK(clknet_leaf_129_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[18]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_013_ ),
    .Q(\i_ibex/id_stage_i/zimm_rs1_type [3]),
    .Q_N(\i_ibex/if_stage_i/_425_ ),
    .CLK(clknet_leaf_135_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[19]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_014_ ),
    .Q(\i_ibex/id_stage_i/zimm_rs1_type [4]),
    .Q_N(\i_ibex/if_stage_i/_424_ ),
    .CLK(clknet_leaf_109_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[1]_reg  (.RESET_B(net1665),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_015_ ),
    .Q(\i_ibex/instr_rdata_id [1]),
    .Q_N(\i_ibex/if_stage_i/_423_ ),
    .CLK(clknet_leaf_107_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[20]_reg  (.CLK(clknet_leaf_129_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_016_ ),
    .Q_N(\i_ibex/if_stage_i/_422_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[21]_reg  (.CLK(clknet_leaf_129_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_017_ ),
    .Q_N(\i_ibex/if_stage_i/_421_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[22]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_018_ ),
    .Q_N(\i_ibex/if_stage_i/_420_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[23]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_019_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [23]),
    .Q_N(\i_ibex/if_stage_i/_419_ ),
    .CLK(clknet_leaf_129_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[24]_reg  (.RESET_B(net1666),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_020_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [24]),
    .Q_N(\i_ibex/if_stage_i/_418_ ),
    .CLK(clknet_leaf_107_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[25]_reg  (.CLK(clknet_leaf_106_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_021_ ),
    .Q_N(\i_ibex/if_stage_i/_417_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[26]_reg  (.CLK(clknet_leaf_107_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_022_ ),
    .Q_N(\i_ibex/if_stage_i/_416_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[27]_reg  (.CLK(clknet_leaf_106_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_023_ ),
    .Q_N(\i_ibex/if_stage_i/_415_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[28]_reg  (.CLK(clknet_leaf_107_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_024_ ),
    .Q_N(\i_ibex/if_stage_i/_414_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[29]_reg  (.CLK(clknet_leaf_107_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_025_ ),
    .Q_N(\i_ibex/if_stage_i/_413_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[2]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_026_ ),
    .Q_N(\i_ibex/if_stage_i/_412_ ),
    .Q(\i_ibex/instr_rdata_id [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[30]_reg  (.CLK(clknet_leaf_106_clk_i_regs),
    .RESET_B(net1668),
    .D(\i_ibex/if_stage_i/_027_ ),
    .Q_N(\i_ibex/if_stage_i/_411_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[31]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_028_ ),
    .Q_N(\i_ibex/if_stage_i/_410_ ),
    .Q(\i_ibex/id_stage_i/imm_u_type [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[3]_reg  (.CLK(clknet_leaf_112_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_029_ ),
    .Q_N(\i_ibex/if_stage_i/_409_ ),
    .Q(\i_ibex/instr_rdata_id [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[4]_reg  (.CLK(clknet_leaf_105_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_030_ ),
    .Q_N(\i_ibex/if_stage_i/_408_ ),
    .Q(\i_ibex/instr_rdata_id [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[5]_reg  (.CLK(clknet_leaf_105_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_031_ ),
    .Q_N(\i_ibex/if_stage_i/_407_ ),
    .Q(\i_ibex/instr_rdata_id [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_alu_id_o[6]_reg  (.CLK(clknet_leaf_105_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_032_ ),
    .Q_N(\i_ibex/if_stage_i/_406_ ),
    .Q(\i_ibex/instr_rdata_id [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[7]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_033_ ),
    .Q(\i_ibex/id_stage_i/imm_s_type [0]),
    .Q_N(\i_ibex/if_stage_i/_405_ ),
    .CLK(clknet_leaf_128_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[8]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_034_ ),
    .Q(\i_ibex/id_stage_i/imm_s_type [1]),
    .Q_N(\i_ibex/if_stage_i/_404_ ),
    .CLK(clknet_leaf_129_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/instr_rdata_alu_id_o[9]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_035_ ),
    .Q(\i_ibex/id_stage_i/imm_s_type [2]),
    .Q_N(\i_ibex/if_stage_i/_403_ ),
    .CLK(clknet_leaf_128_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[0]_reg  (.CLK(clknet_leaf_110_clk_i_regs),
    .RESET_B(net1668),
    .D(\i_ibex/if_stage_i/_036_ ),
    .Q_N(\i_ibex/if_stage_i/_402_ ),
    .Q(\i_ibex/instr_rdata_c_id [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[10]_reg  (.CLK(clknet_leaf_109_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_037_ ),
    .Q_N(\i_ibex/if_stage_i/_401_ ),
    .Q(\i_ibex/instr_rdata_c_id [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[11]_reg  (.CLK(clknet_5_17__leaf_clk_i_regs),
    .RESET_B(net1668),
    .D(\i_ibex/if_stage_i/_038_ ),
    .Q_N(\i_ibex/if_stage_i/_400_ ),
    .Q(\i_ibex/instr_rdata_c_id [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[12]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_039_ ),
    .Q_N(\i_ibex/if_stage_i/_399_ ),
    .Q(\i_ibex/instr_rdata_c_id [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[13]_reg  (.CLK(clknet_leaf_109_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_040_ ),
    .Q_N(\i_ibex/if_stage_i/_398_ ),
    .Q(\i_ibex/instr_rdata_c_id [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[14]_reg  (.CLK(clknet_5_17__leaf_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_041_ ),
    .Q_N(\i_ibex/if_stage_i/_397_ ),
    .Q(\i_ibex/instr_rdata_c_id [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[15]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_042_ ),
    .Q_N(\i_ibex/if_stage_i/_396_ ),
    .Q(\i_ibex/instr_rdata_c_id [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[1]_reg  (.CLK(clknet_leaf_110_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_043_ ),
    .Q_N(\i_ibex/if_stage_i/_395_ ),
    .Q(\i_ibex/instr_rdata_c_id [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[2]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_044_ ),
    .Q_N(\i_ibex/if_stage_i/_394_ ),
    .Q(\i_ibex/instr_rdata_c_id [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[3]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/_045_ ),
    .Q_N(\i_ibex/if_stage_i/_393_ ),
    .Q(\i_ibex/instr_rdata_c_id [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[4]_reg  (.CLK(clknet_leaf_108_clk_i_regs),
    .RESET_B(net1666),
    .D(\i_ibex/if_stage_i/_046_ ),
    .Q_N(\i_ibex/if_stage_i/_392_ ),
    .Q(\i_ibex/instr_rdata_c_id [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[5]_reg  (.CLK(clknet_leaf_107_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_047_ ),
    .Q_N(\i_ibex/if_stage_i/_391_ ),
    .Q(\i_ibex/instr_rdata_c_id [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[6]_reg  (.CLK(clknet_leaf_107_clk_i_regs),
    .RESET_B(net1667),
    .D(\i_ibex/if_stage_i/_048_ ),
    .Q_N(\i_ibex/if_stage_i/_390_ ),
    .Q(\i_ibex/instr_rdata_c_id [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[7]_reg  (.CLK(clknet_leaf_109_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_049_ ),
    .Q_N(\i_ibex/if_stage_i/_389_ ),
    .Q(\i_ibex/instr_rdata_c_id [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[8]_reg  (.CLK(clknet_leaf_109_clk_i_regs),
    .RESET_B(net1668),
    .D(\i_ibex/if_stage_i/_050_ ),
    .Q_N(\i_ibex/if_stage_i/_388_ ),
    .Q(\i_ibex/instr_rdata_c_id [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_rdata_c_id_o[9]_reg  (.CLK(clknet_leaf_109_clk_i_regs),
    .RESET_B(net1665),
    .D(\i_ibex/if_stage_i/_051_ ),
    .Q_N(\i_ibex/if_stage_i/_440_ ),
    .Q(\i_ibex/instr_rdata_c_id [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/instr_valid_id_o_reg  (.CLK(clknet_leaf_89_clk_i_regs),
    .RESET_B(net1576),
    .D(\i_ibex/if_stage_i/instr_valid_id_d ),
    .Q_N(\i_ibex/if_stage_i/_387_ ),
    .Q(\i_ibex/instr_valid_id ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[0]_reg  (.RESET_B(net1576),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_052_ ),
    .Q(\i_ibex/pc_id [0]),
    .Q_N(\i_ibex/if_stage_i/_386_ ),
    .CLK(clknet_leaf_83_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[10]_reg  (.RESET_B(net1533),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_053_ ),
    .Q(\i_ibex/pc_id [10]),
    .Q_N(\i_ibex/if_stage_i/_385_ ),
    .CLK(clknet_leaf_95_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[11]_reg  (.RESET_B(net1533),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_054_ ),
    .Q(\i_ibex/pc_id [11]),
    .Q_N(\i_ibex/if_stage_i/_384_ ),
    .CLK(clknet_leaf_95_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[12]_reg  (.RESET_B(net1567),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_055_ ),
    .Q(\i_ibex/pc_id [12]),
    .Q_N(\i_ibex/if_stage_i/_383_ ),
    .CLK(clknet_leaf_95_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[13]_reg  (.RESET_B(net1594),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_056_ ),
    .Q(\i_ibex/pc_id [13]),
    .Q_N(\i_ibex/if_stage_i/_382_ ),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[14]_reg  (.RESET_B(net1567),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_057_ ),
    .Q(\i_ibex/pc_id [14]),
    .Q_N(\i_ibex/if_stage_i/_381_ ),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[15]_reg  (.RESET_B(net1594),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_058_ ),
    .Q(\i_ibex/pc_id [15]),
    .Q_N(\i_ibex/if_stage_i/_380_ ),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[16]_reg  (.RESET_B(net1596),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_059_ ),
    .Q(\i_ibex/pc_id [16]),
    .Q_N(\i_ibex/if_stage_i/_379_ ),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[17]_reg  (.RESET_B(net1596),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_060_ ),
    .Q(\i_ibex/pc_id [17]),
    .Q_N(\i_ibex/if_stage_i/_378_ ),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[18]_reg  (.RESET_B(net1634),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_061_ ),
    .Q(\i_ibex/pc_id [18]),
    .Q_N(\i_ibex/if_stage_i/_377_ ),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[19]_reg  (.RESET_B(net1633),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_062_ ),
    .Q(\i_ibex/pc_id [19]),
    .Q_N(\i_ibex/if_stage_i/_376_ ),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[1]_reg  (.RESET_B(net1549),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_063_ ),
    .Q(\i_ibex/pc_id [1]),
    .Q_N(\i_ibex/if_stage_i/_375_ ),
    .CLK(clknet_leaf_83_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[20]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_064_ ),
    .Q(\i_ibex/pc_id [20]),
    .Q_N(\i_ibex/if_stage_i/_374_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[21]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_065_ ),
    .Q(\i_ibex/pc_id [21]),
    .Q_N(\i_ibex/if_stage_i/_373_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[22]_reg  (.RESET_B(net1626),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_066_ ),
    .Q(\i_ibex/pc_id [22]),
    .Q_N(\i_ibex/if_stage_i/_372_ ),
    .CLK(clknet_leaf_138_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[23]_reg  (.RESET_B(net1628),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_067_ ),
    .Q(\i_ibex/pc_id [23]),
    .Q_N(\i_ibex/if_stage_i/_371_ ),
    .CLK(clknet_leaf_137_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[24]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_068_ ),
    .Q(\i_ibex/pc_id [24]),
    .Q_N(\i_ibex/if_stage_i/_370_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[25]_reg  (.RESET_B(net1628),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_069_ ),
    .Q(\i_ibex/pc_id [25]),
    .Q_N(\i_ibex/if_stage_i/_369_ ),
    .CLK(clknet_leaf_137_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[26]_reg  (.RESET_B(net1596),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_070_ ),
    .Q(\i_ibex/pc_id [26]),
    .Q_N(\i_ibex/if_stage_i/_368_ ),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[27]_reg  (.RESET_B(net1592),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_071_ ),
    .Q(\i_ibex/pc_id [27]),
    .Q_N(\i_ibex/if_stage_i/_367_ ),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[28]_reg  (.RESET_B(net1592),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_072_ ),
    .Q(\i_ibex/pc_id [28]),
    .Q_N(\i_ibex/if_stage_i/_366_ ),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[29]_reg  (.RESET_B(net1593),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_073_ ),
    .Q(\i_ibex/pc_id [29]),
    .Q_N(\i_ibex/if_stage_i/_365_ ),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[2]_reg  (.RESET_B(net1549),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_074_ ),
    .Q(\i_ibex/pc_id [2]),
    .Q_N(\i_ibex/if_stage_i/_364_ ),
    .CLK(clknet_leaf_82_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[30]_reg  (.RESET_B(net1633),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_075_ ),
    .Q(\i_ibex/pc_id [30]),
    .Q_N(\i_ibex/if_stage_i/_363_ ),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[31]_reg  (.RESET_B(net1596),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_076_ ),
    .Q(\i_ibex/pc_id [31]),
    .Q_N(\i_ibex/if_stage_i/_362_ ),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[3]_reg  (.RESET_B(net1575),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_077_ ),
    .Q(\i_ibex/pc_id [3]),
    .Q_N(\i_ibex/if_stage_i/_361_ ),
    .CLK(clknet_leaf_82_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[4]_reg  (.RESET_B(net1546),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_078_ ),
    .Q(\i_ibex/pc_id [4]),
    .Q_N(\i_ibex/if_stage_i/_360_ ),
    .CLK(clknet_leaf_92_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[5]_reg  (.RESET_B(net1575),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_079_ ),
    .Q(\i_ibex/pc_id [5]),
    .Q_N(\i_ibex/if_stage_i/_359_ ),
    .CLK(clknet_leaf_92_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[6]_reg  (.RESET_B(net1575),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_080_ ),
    .Q(\i_ibex/pc_id [6]),
    .Q_N(\i_ibex/if_stage_i/_358_ ),
    .CLK(clknet_leaf_92_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[7]_reg  (.RESET_B(net1575),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_081_ ),
    .Q(\i_ibex/pc_id [7]),
    .Q_N(\i_ibex/if_stage_i/_357_ ),
    .CLK(clknet_leaf_93_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[8]_reg  (.RESET_B(net1567),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_082_ ),
    .Q(\i_ibex/pc_id [8]),
    .Q_N(\i_ibex/if_stage_i/_356_ ),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/pc_id_o[9]_reg  (.RESET_B(net1533),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/_083_ ),
    .Q(\i_ibex/pc_id [9]),
    .Q_N(\i_ibex/if_stage_i/_355_ ),
    .CLK(clknet_leaf_95_clk_i_regs));
 sg13g2_buf_8 fanout499 (.A(net517),
    .X(net499),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(net517),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(net517),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout496 (.A(net515),
    .X(net496),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(\i_ibex/cs_registers_i/_0873_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(net495),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_424_  (.B1(net1466),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_066_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/discard_req_q ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_425_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_067_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [0]),
    .B(net1673),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout493 (.A(net495),
    .X(net493),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(net495),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_428_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1120),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [1]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_070_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q [1]));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_429_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_070_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_071_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_066_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_067_ ));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_430_  (.A(net1671),
    .B_N(\i_ibex/if_stage_i/prefetch_buffer_i/_071_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_s [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_431_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_072_ ),
    .A(net1673),
    .VSS(VSS));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net495),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_433_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1120),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [0]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_074_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q [0]));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_434_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_074_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_075_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_072_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_066_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_435_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_075_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_071_ ),
    .S(net1671),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_s [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_436_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_076_ ),
    .A(net1124),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_437_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_077_ ),
    .B(net698),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [1]));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_438_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_078_ ),
    .B(net1484),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [0]));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_439_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_077_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_078_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_440_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_080_ ),
    .A(net475),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_441_  (.A(\i_ibex/instr_req_gated ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__Y_B ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/if_stage_i/prefetch_buffer_i/_442_  (.A2(\i_ibex/if_stage_i/prefetch_buffer_i/_081_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_080_ ),
    .B1(net1466),
    .X(instr_req_o),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_443_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [0]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [1]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_444_  (.Y(\i_ibex/if_busy ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_082_ ),
    .A_N(instr_req_o),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_445_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/discard_req_d ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_066_ ),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_446_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__A_B ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__Y_B ),
    .A(\i_ibex/instr_req_gated ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_083_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/if_stage_i/prefetch_buffer_i/_447_  (.A(net1125),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_079_ ),
    .C(net1321),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(\i_ibex/alu_operand_b_ex [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_449_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_086_ ),
    .B1(net1030),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [10]),
    .A2(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .A1(net1123),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_450_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_087_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_086_ ),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_451_  (.A(\i_ibex/if_stage_i/fetch_addr_n [3]),
    .B(\i_ibex/if_stage_i/fetch_addr_n [2]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_452_  (.B(\i_ibex/if_stage_i/fetch_addr_n [5]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [4]),
    .A(net1118),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_089_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_088_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_453_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_090_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [3]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_454_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_077_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_078_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_091_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_090_ ));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_455_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [5]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [4]),
    .A(net475),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_091_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_456_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_093_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [9]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_457_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_094_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [6]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_458_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_095_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [8]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_459_  (.A(net1118),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_093_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_094_ ),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_095_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_096_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_460_  (.A(\i_ibex/if_stage_i/fetch_addr_n [8]),
    .B(\i_ibex/if_stage_i/fetch_addr_n [7]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_461_  (.B(\i_ibex/if_stage_i/fetch_addr_n [9]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [6]),
    .A(net1118),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_098_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_097_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_462_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_098_ ),
    .C1(net1321),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_096_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_089_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_099_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_092_ ));
 sg13g2_buf_8 fanout489 (.A(net490),
    .X(net489),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/prefetch_buffer_i/_464_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1321),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_078_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_077_ ));
 sg13g2_nor2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_465_  (.A(net1125),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net489),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_467_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_104_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [10]),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_468_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [10]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_469_  (.A(net411),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_105_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_470_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_104_ ),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_106_ ),
    .B1(net1029),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_087_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_000_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_099_ ));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net489),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_472_  (.A(\i_ibex/if_stage_i/fetch_addr_n [11]),
    .B_N(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_473_  (.A(net1124),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [11]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_104_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_109_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_474_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1118),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_108_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_110_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_109_ ));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/prefetch_buffer_i/_475_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1321),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_111_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_092_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_089_ ));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/prefetch_buffer_i/_476_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1029),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_112_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_098_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_096_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_477_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_113_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_111_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout486 (.A(net489),
    .X(net486),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_479_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [11]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [11]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_480_  (.A(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .B_N(\i_ibex/if_stage_i/fetch_addr_n [11]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 max_cap485 (.A(net1099),
    .X(net485),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(\i_ibex/csr_addr [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout483 (.A(\i_ibex/csr_addr [5]),
    .X(net483),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_484_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/_120_ ),
    .A(net475),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [11]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_485_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1124),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_120_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_116_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_113_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_121_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_115_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_486_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_121_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_001_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_110_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_113_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_487_  (.B(\i_ibex/if_stage_i/fetch_addr_n [11]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .A(net1116),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_488_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [11]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [10]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_123_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1123));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_489_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_124_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_122_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_490_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_125_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_099_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_491_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_126_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [12]),
    .VSS(VSS));
 sg13g2_and2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_492_  (.A(net475),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout482 (.A(\i_ibex/cs_registers_i/_0942_ ),
    .X(net482),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_494_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_129_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [12]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_495_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_130_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_129_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_126_ ),
    .A1(net1123),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout481 (.A(\i_ibex/cs_registers_i/_0942_ ),
    .X(net481),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_497_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_132_ ),
    .A(net1116),
    .B(\i_ibex/if_stage_i/fetch_addr_n [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_498_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_132_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_133_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_129_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_499_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_134_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_125_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_133_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_102_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_500_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_134_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_002_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_125_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_130_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_501_  (.B(\i_ibex/if_stage_i/fetch_addr_n [13]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_126_ ),
    .A(net1117),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_502_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_136_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [12]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_503_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [13]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_136_ ),
    .A(net476),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_504_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [13]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_129_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_138_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_505_  (.A(\i_ibex/if_stage_i/fetch_addr_n [13]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_132_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_139_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_506_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1030),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_138_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_140_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_139_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_507_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_137_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_140_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_135_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_508_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [13]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [13]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_509_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_141_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_142_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/_125_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_510_  (.B(\i_ibex/if_stage_i/fetch_addr_n [13]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [12]),
    .A(net1116),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_143_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_511_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [13]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [12]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_144_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net1123));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_512_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_145_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_143_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_144_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_123_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_513_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_146_ ),
    .A(net411),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_514_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_147_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [14]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_515_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_148_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [14]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_516_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_149_ ),
    .B1(net1030),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_148_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_147_ ),
    .A1(net1123),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_517_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_150_ ),
    .A(net1116),
    .B(\i_ibex/if_stage_i/fetch_addr_n [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_518_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_150_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_151_ ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_148_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_519_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_152_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_146_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_151_ ),
    .A2(net1028),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_520_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_152_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_004_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_146_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_149_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_521_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_153_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [14]),
    .B(net1030),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_522_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_150_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_153_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_154_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_146_ ));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_523_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [15]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [15]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_524_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_155_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_154_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_525_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [16]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [16]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_156_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_526_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_157_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [15]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_527_  (.B(\i_ibex/if_stage_i/fetch_addr_n [15]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [14]),
    .A(net1116),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_528_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_158_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_159_ ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_157_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_529_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_159_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_160_ ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_530_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_146_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_160_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_531_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_161_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_156_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_532_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_162_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [17]),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_533_  (.A(net411),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_145_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_156_ ),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_159_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_534_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_164_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [17]),
    .A2(\i_ibex/if_stage_i/fetch_addr_n [17]),
    .A1(net1123),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_535_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_165_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_164_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_536_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [17]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [17]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_166_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_537_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_163_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_166_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_538_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_165_ ),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_167_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_163_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_162_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_007_ ),
    .A2(net1028));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_539_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_168_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [17]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_540_  (.B(\i_ibex/if_stage_i/fetch_addr_n [17]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [16]),
    .A(net1117),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_541_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_169_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_170_ ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_168_ ));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_542_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/_171_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_145_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_159_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_170_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_543_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_112_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_171_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_111_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_172_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_544_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_173_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [18]),
    .VSS(VSS));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_546_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_175_ ),
    .A(net1119),
    .B(\i_ibex/if_stage_i/fetch_addr_n [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_547_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_175_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_176_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_173_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_548_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_008_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_172_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_549_  (.A(\i_ibex/if_stage_i/fetch_addr_n [19]),
    .B_N(\i_ibex/if_stage_i/fetch_addr_n [18]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_177_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_550_  (.A(net1124),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [19]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_173_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_551_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1119),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_177_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_179_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_178_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_552_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [19]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [19]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_180_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_553_  (.A(\i_ibex/if_stage_i/fetch_addr_n [18]),
    .B_N(\i_ibex/if_stage_i/fetch_addr_n [19]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_181_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_554_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/_182_ ),
    .A(net475),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [19]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_173_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_555_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1124),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_182_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_181_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_172_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_183_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_180_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_556_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_183_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_009_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_172_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_179_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_557_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_184_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [19]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_558_  (.B(\i_ibex/if_stage_i/fetch_addr_n [19]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [18]),
    .A(net1117),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_559_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_185_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_186_ ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_184_ ));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_560_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_159_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_170_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_145_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_187_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_186_ ));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_561_  (.A(net1028),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_187_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_562_  (.A(net411),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_188_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_563_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [20]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [20]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_564_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_190_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_189_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_565_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_191_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [20]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_566_  (.B(\i_ibex/if_stage_i/fetch_addr_n [20]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [21]),
    .A(net1114),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_567_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_192_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_193_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_191_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_568_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [21]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [21]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_569_  (.A(\i_ibex/if_stage_i/fetch_addr_n [20]),
    .B(\i_ibex/if_stage_i/fetch_addr_n [21]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_195_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_570_  (.A(net1122),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [20]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [21]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_571_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1114),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_195_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_197_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_196_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_572_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_197_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_198_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_189_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_194_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_573_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_189_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_193_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_011_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_198_ ));
 sg13g2_nor2b_2 \i_ibex/if_stage_i/prefetch_buffer_i/_574_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_187_ ),
    .B_N(\i_ibex/if_stage_i/prefetch_buffer_i/_193_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_199_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_575_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_112_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_199_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_111_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_576_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_201_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [22]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_577_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_202_ ),
    .A(net1116),
    .B(\i_ibex/if_stage_i/fetch_addr_n [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_578_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_202_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_203_ ),
    .VSS(VSS),
    .A1(net1129),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_201_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_579_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_012_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_200_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_203_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_580_  (.A(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .B_N(\i_ibex/if_stage_i/fetch_addr_n [22]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_581_  (.A(net1123),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [23]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_201_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_582_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1116),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_204_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_206_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_205_ ));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_583_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [23]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .S(net1139),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_584_  (.A(\i_ibex/if_stage_i/fetch_addr_n [22]),
    .B_N(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_208_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_585_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/_209_ ),
    .A(net475),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [23]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_201_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_586_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1123),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_209_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_208_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_200_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_210_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_207_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_587_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_210_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_013_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_200_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_206_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_588_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_211_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [23]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_589_  (.B(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [22]),
    .A(net1117),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_212_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_590_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_212_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_213_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_211_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_591_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_199_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_213_ ),
    .A(net411),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_214_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_592_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_215_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [24]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_593_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_216_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [24]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_594_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_217_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_216_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_215_ ),
    .A1(net1122),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_595_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_218_ ),
    .A(net1114),
    .B(\i_ibex/if_stage_i/fetch_addr_n [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_596_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_218_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_219_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_216_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_597_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_220_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_214_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_219_ ),
    .A2(net1028),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_598_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_220_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_014_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_214_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_217_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_599_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_221_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [24]),
    .B(net1030),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_600_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_218_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_221_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_222_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_214_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_601_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [25]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [25]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_223_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_602_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_223_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_222_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_603_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_224_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [25]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_604_  (.B(\i_ibex/if_stage_i/fetch_addr_n [25]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [24]),
    .A(net1114),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_225_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_605_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_225_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_226_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_224_ ));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_606_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_199_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_213_ ),
    .A(net411),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_226_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_607_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_228_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [26]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_608_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_229_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [26]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_609_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_230_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_229_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_228_ ),
    .A1(net1122),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_610_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_231_ ),
    .A(net1114),
    .B(\i_ibex/if_stage_i/fetch_addr_n [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_611_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_231_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_232_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_229_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_612_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_233_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_227_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_232_ ),
    .A2(net1028),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_613_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_233_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_016_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_227_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_230_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_614_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_234_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [27]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_615_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_235_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [27]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_616_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_236_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_235_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_234_ ),
    .A1(net1122),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_617_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [25]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [24]),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [26]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_618_  (.B(\i_ibex/if_stage_i/fetch_addr_n [26]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [25]),
    .A(net1114),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_238_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/fetch_addr_n [24]));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_619_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_238_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_239_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_237_ ));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_620_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_199_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_213_ ),
    .A(net411),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_240_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_239_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_621_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_241_ ),
    .A(net1114),
    .B(\i_ibex/if_stage_i/fetch_addr_n [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_622_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_241_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_242_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_235_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_623_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_243_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_240_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_242_ ),
    .A2(net1028),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_624_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_243_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_017_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_236_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_240_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_625_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [23]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [22]),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [27]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_626_  (.B(\i_ibex/if_stage_i/fetch_addr_n [27]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .A(net1117),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_245_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/fetch_addr_n [22]));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_627_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_245_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_246_ ),
    .VSS(VSS),
    .A1(net1127),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_244_ ));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_628_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_199_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_239_ ),
    .A(net411),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_247_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_246_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_629_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_248_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [28]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_630_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_249_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [28]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_631_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_250_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_249_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_248_ ),
    .A1(net1122),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_632_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_251_ ),
    .A(net1114),
    .B(\i_ibex/if_stage_i/fetch_addr_n [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_633_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_251_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_252_ ),
    .VSS(VSS),
    .A1(net1128),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_249_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_634_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_253_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_247_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_252_ ),
    .A2(net1028),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_635_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_253_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_018_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_247_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_250_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_636_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_254_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [28]),
    .B(net1030),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_637_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_251_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_254_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_255_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_247_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_638_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [29]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [29]),
    .S(net1139),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_256_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_639_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_256_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_255_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_640_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_257_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [2]),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_641_  (.A(net1125),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_079_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_642_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_259_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [2]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_643_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_260_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_258_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_259_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_257_ ),
    .A1(net1125),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_644_  (.A(net1125),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_259_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_261_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_645_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_262_ ),
    .A(net1120),
    .B(\i_ibex/if_stage_i/fetch_addr_n [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_646_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_262_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_263_ ),
    .VSS(VSS),
    .A1(net1131),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_259_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_647_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_264_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_263_ ),
    .B2(net1321),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_261_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_648_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_264_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_020_ ),
    .VSS(VSS),
    .A1(net1321),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_260_ ));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_649_  (.B(\i_ibex/if_stage_i/fetch_addr_n [29]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [28]),
    .A(net1115),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_265_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_650_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [29]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [28]),
    .A(net476),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_651_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_265_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_266_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_267_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_247_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_652_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [30]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [30]),
    .S(net1139),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_653_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_268_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_267_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_654_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_269_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [31]),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_655_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [30]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [29]),
    .A(net476),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_270_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [28]));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_656_  (.B(\i_ibex/if_stage_i/fetch_addr_n [30]),
    .C(\i_ibex/if_stage_i/fetch_addr_n [29]),
    .A(net1115),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_271_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/fetch_addr_n [28]));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_657_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_270_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_271_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_272_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_658_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_273_ ),
    .B(net1115),
    .A_N(\i_ibex/if_stage_i/fetch_addr_n [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_659_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_273_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_274_ ),
    .VSS(VSS),
    .A1(net1128),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [31]));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_660_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_275_ ),
    .A(net1115),
    .B(\i_ibex/if_stage_i/fetch_addr_n [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_661_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_276_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [31]),
    .B(net1030),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_662_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_275_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_276_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_277_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_272_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_663_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_274_ ),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_277_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_272_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_269_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_278_ ),
    .A2(net1028));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_664_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_275_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_279_ ),
    .VSS(VSS),
    .A1(net1128),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_269_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_665_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_278_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_279_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/_247_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_666_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_280_ ),
    .A(net1120),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_667_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_281_ ),
    .A(net476),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_091_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_668_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_280_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_281_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_282_ ),
    .B1(net1321));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_669_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_258_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_283_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [3]),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [2]));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_670_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_262_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_283_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_284_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_083_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_671_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1120),
    .A2(\i_ibex/if_stage_i/fetch_addr_n [3]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_285_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_284_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_672_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_286_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [3]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_673_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_286_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_023_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_282_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_285_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_674_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_287_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_282_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_675_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_288_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [4]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_676_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_289_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [4]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_677_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_290_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_084_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_289_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_288_ ),
    .A1(net1124),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_678_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_291_ ),
    .A(net1121),
    .B(\i_ibex/if_stage_i/fetch_addr_n [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_679_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_291_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_292_ ),
    .VSS(VSS),
    .A1(net1131),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_289_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_680_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_293_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_287_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_292_ ),
    .A2(net1029),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_681_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_293_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_024_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_287_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_290_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_682_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_294_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [5]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_683_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_295_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_282_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_292_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_684_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_296_ ),
    .B(net1120),
    .A_N(\i_ibex/if_stage_i/fetch_addr_n [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_685_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_296_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_297_ ),
    .VSS(VSS),
    .A1(net1131),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [5]));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_686_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_298_ ),
    .A(net1121),
    .B(\i_ibex/if_stage_i/fetch_addr_n [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_687_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_299_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [5]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_688_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_298_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_299_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_300_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_295_ ));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_689_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_297_ ),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/_300_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_295_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_294_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_025_ ),
    .A2(net1029));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_690_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_301_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_111_ ),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_691_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_302_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [6]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_692_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_303_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_084_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_094_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_302_ ),
    .A1(net1124),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_693_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_304_ ),
    .A(net1118),
    .B(\i_ibex/if_stage_i/fetch_addr_n [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_694_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_305_ ),
    .A(net476),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_695_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_306_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_304_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_696_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_307_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_306_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_301_ ),
    .A2(net1029),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_697_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_307_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_026_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_301_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_303_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_698_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_308_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_111_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_306_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_699_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_309_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [7]),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_700_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_310_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [7]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_701_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_311_ ),
    .B1(net1030),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_310_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_309_ ),
    .A1(net1124),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_702_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_312_ ),
    .A(net1119),
    .B(\i_ibex/if_stage_i/fetch_addr_n [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_703_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_312_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_313_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_310_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_704_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_314_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_308_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_313_ ),
    .A2(net1029),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_705_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_314_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_027_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_308_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_311_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_706_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_315_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [8]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_707_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_316_ ),
    .A(net1119),
    .B(\i_ibex/if_stage_i/fetch_addr_n [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_708_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_316_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_317_ ),
    .VSS(VSS),
    .A1(net1131),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_315_ ));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_709_  (.A(net475),
    .B(\i_ibex/if_stage_i/fetch_addr_n [8]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_309_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_318_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/_710_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/_315_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [7]),
    .A(net476),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_711_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_320_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_319_ ),
    .A_N(\i_ibex/if_stage_i/prefetch_buffer_i/_318_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_712_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_305_ ),
    .C1(net1321),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_304_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_089_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_321_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_092_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_713_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_317_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_320_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/_321_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_714_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [7]),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_323_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_315_ ));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_715_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_324_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_101_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [8]));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_716_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_324_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_325_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_322_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_323_ ));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_717_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [8]),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_309_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_326_ ),
    .B1(net475));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_718_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_322_ ),
    .B_N(\i_ibex/if_stage_i/prefetch_buffer_i/_326_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_327_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_719_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net476),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_325_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_028_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_327_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_720_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_328_ ),
    .A(net1118),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_721_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_328_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_329_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_095_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_722_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_330_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_321_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/_329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_723_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_331_ ),
    .A(\i_ibex/if_stage_i/fetch_addr_n [9]),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_724_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_332_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_127_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_093_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_331_ ),
    .A1(net1125),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_725_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_333_ ),
    .A(net1118),
    .B(\i_ibex/if_stage_i/fetch_addr_n [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_726_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_333_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_334_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_093_ ));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_727_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_335_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_330_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_334_ ),
    .A2(net1029),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_728_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_335_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_029_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_330_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_332_ ));
 sg13g2_and2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_729_  (.A(net1671),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid_$_AND__Y_B ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net481),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_731_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_279_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [31]),
    .S(net1467),
    .X(instr_addr_o[31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_732_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_268_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [30]),
    .S(net1466),
    .X(instr_addr_o[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_733_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_194_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [21]),
    .S(net1465),
    .X(instr_addr_o[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_734_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_190_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [20]),
    .S(net1467),
    .X(instr_addr_o[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_735_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_180_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [19]),
    .S(net1466),
    .X(instr_addr_o[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_736_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_176_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [18]),
    .S(net1469),
    .X(instr_addr_o[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_737_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_337_ ),
    .A(net1116),
    .B(\i_ibex/if_stage_i/fetch_addr_n [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_738_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_337_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_338_ ),
    .VSS(VSS),
    .A1(net1132),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_162_ ));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_739_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_338_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [17]),
    .S(net1465),
    .X(instr_addr_o[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_740_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_156_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [16]),
    .S(net1466),
    .X(instr_addr_o[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_741_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_155_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [15]),
    .S(net1467),
    .X(instr_addr_o[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_742_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_151_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [14]),
    .S(net1467),
    .X(instr_addr_o[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(net481),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_744_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_142_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [13]),
    .S(net1465),
    .X(instr_addr_o[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_745_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_133_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [12]),
    .S(net1467),
    .X(instr_addr_o[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_746_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_256_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [29]),
    .S(net1465),
    .X(instr_addr_o[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_747_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_115_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [11]),
    .S(net1469),
    .X(instr_addr_o[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_748_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_340_ ),
    .A(net1118),
    .B(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_749_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_340_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_341_ ),
    .VSS(VSS),
    .A1(net1130),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_104_ ));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_750_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_341_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [10]),
    .S(net1468),
    .X(instr_addr_o[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_751_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_334_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [9]),
    .S(net1468),
    .X(instr_addr_o[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_752_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_317_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [8]),
    .S(net1468),
    .X(instr_addr_o[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_753_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_313_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [7]),
    .S(net1465),
    .X(instr_addr_o[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_754_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_306_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [6]),
    .S(net1465),
    .X(instr_addr_o[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_755_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_298_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_342_ ),
    .VSS(VSS),
    .A1(net1131),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_294_ ));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_756_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_342_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [5]),
    .S(net1467),
    .X(instr_addr_o[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(net481),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_758_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_292_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [4]),
    .S(net1467),
    .X(instr_addr_o[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_759_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [3]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [3]),
    .S(net1138),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_344_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_760_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_344_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [3]),
    .S(net1466),
    .X(instr_addr_o[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_761_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_263_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [2]),
    .S(net1467),
    .X(instr_addr_o[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_762_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_252_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [28]),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/valid_req_q ),
    .X(instr_addr_o[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_763_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_242_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [27]),
    .S(net1468),
    .X(instr_addr_o[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_764_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_232_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [26]),
    .S(net1465),
    .X(instr_addr_o[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_765_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_223_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [25]),
    .S(net1465),
    .X(instr_addr_o[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_766_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_219_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [24]),
    .S(net1468),
    .X(instr_addr_o[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_767_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_207_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [23]),
    .S(net1468),
    .X(instr_addr_o[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/_768_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/_203_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [22]),
    .S(net1466),
    .X(instr_addr_o[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/_769_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_345_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [1]),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/_770_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_346_ ),
    .B(instr_req_o),
    .A_N(\i_ibex/if_stage_i/prefetch_buffer_i/_067_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_771_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/_345_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_346_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_s [1]),
    .B1(net1671));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_772_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_347_ ),
    .A(net1673),
    .B(instr_req_o),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_773_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/_348_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_345_ ),
    .B(net1671),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/_774_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/_348_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_349_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [0]),
    .A2(net1671));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/_775_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_s [0]),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/_347_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/_349_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/_082_ ),
    .A1(net1671),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/_776_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__A_B ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/_080_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/_072_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/_350_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_081_ ));
 sg13g2_buf_2 fanout476 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_076_ ),
    .X(net476),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_778_  (.A0(instr_addr_o[10]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [10]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_779_  (.A0(instr_addr_o[11]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [11]),
    .S(net1027),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_780_  (.A0(instr_addr_o[12]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [12]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_781_  (.A0(instr_addr_o[13]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [13]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_782_  (.A0(instr_addr_o[14]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [14]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_783_  (.A0(instr_addr_o[15]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [15]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_784_  (.A0(instr_addr_o[16]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [16]),
    .S(net1024),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_785_  (.A0(instr_addr_o[17]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [17]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_786_  (.A0(instr_addr_o[18]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [18]),
    .S(net1027),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_787_  (.A0(instr_addr_o[19]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [19]),
    .S(net1024),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout475 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_076_ ),
    .X(net475),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_789_  (.A0(instr_addr_o[20]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [20]),
    .S(net1026),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_790_  (.A0(instr_addr_o[21]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [21]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_791_  (.A0(instr_addr_o[22]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [22]),
    .S(net1024),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_792_  (.A0(instr_addr_o[23]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [23]),
    .S(net1026),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_793_  (.A0(instr_addr_o[24]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [24]),
    .S(net1026),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_794_  (.A0(instr_addr_o[25]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [25]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_795_  (.A0(instr_addr_o[26]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [26]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_796_  (.A0(instr_addr_o[27]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [27]),
    .S(net1026),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_797_  (.A0(instr_addr_o[28]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [28]),
    .S(net1024),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_798_  (.A0(instr_addr_o[29]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [29]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 max_cap474 (.A(net1057),
    .X(net474),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_800_  (.A0(instr_addr_o[2]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [2]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_801_  (.A0(instr_addr_o[30]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [30]),
    .S(net1024),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_802_  (.A0(instr_addr_o[31]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [31]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_803_  (.A0(instr_addr_o[3]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [3]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_804_  (.A0(instr_addr_o[4]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [4]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_805_  (.A0(instr_addr_o[5]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [5]),
    .S(net1025),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_806_  (.A0(instr_addr_o[6]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [6]),
    .S(net1024),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_807_  (.A0(instr_addr_o[7]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [7]),
    .S(net1023),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_808_  (.A0(instr_addr_o[8]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [8]),
    .S(net1026),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_058_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_809_  (.A0(instr_addr_o[9]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [9]),
    .S(net1026),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/_810_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_072_ ),
    .B(instr_req_o),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/valid_req_d ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \i_ibex/cs_registers_i/_2163__378  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net378));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q[0]_reg  (.CLK(clknet_leaf_142_clk_i_regs),
    .RESET_B(net1562),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_s [0]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid_$_AND__Y_B ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q[1]_reg  (.CLK(clknet_leaf_142_clk_i_regs),
    .RESET_B(net1652),
    .D(net1672),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_413_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/discard_req_q_reg  (.CLK(clknet_leaf_143_clk_i_regs),
    .RESET_B(net1652),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/discard_req_d ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_412_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/discard_req_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[10]_reg  (.CLK(clknet_leaf_150_clk_i_regs),
    .RESET_B(net1561),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_000_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_411_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[11]_reg  (.CLK(clknet_leaf_147_clk_i_regs),
    .RESET_B(net1560),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_001_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_410_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[12]_reg  (.CLK(clknet_leaf_148_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_002_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_409_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[13]_reg  (.CLK(clknet_leaf_149_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_003_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_408_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[14]_reg  (.CLK(clknet_leaf_149_clk_i_regs),
    .RESET_B(net1582),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_004_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_407_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[15]_reg  (.CLK(clknet_leaf_142_clk_i_regs),
    .RESET_B(net1561),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_005_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_406_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[16]_reg  (.CLK(clknet_leaf_149_clk_i_regs),
    .RESET_B(net1582),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_006_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_405_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[17]_reg  (.CLK(clknet_leaf_153_clk_i_regs),
    .RESET_B(net1583),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_007_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_404_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[18]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1643),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_008_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_403_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[19]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1643),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_009_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_402_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[20]_reg  (.CLK(clknet_leaf_4_clk_i_regs),
    .RESET_B(net1645),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_010_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_401_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[21]_reg  (.CLK(clknet_leaf_152_clk_i_regs),
    .RESET_B(net1625),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_011_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_400_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[22]_reg  (.CLK(clknet_leaf_153_clk_i_regs),
    .RESET_B(net1643),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_012_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_399_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[23]_reg  (.RESET_B(net1583),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_013_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [23]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_398_ ),
    .CLK(clknet_leaf_153_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[24]_reg  (.CLK(clknet_leaf_153_clk_i_regs),
    .RESET_B(net1583),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_014_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_397_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[25]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1625),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_015_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_396_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[26]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1643),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_016_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_395_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[27]_reg  (.CLK(clknet_leaf_153_clk_i_regs),
    .RESET_B(net1643),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_017_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_394_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[28]_reg  (.CLK(clknet_leaf_152_clk_i_regs),
    .RESET_B(net1583),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_018_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_393_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[29]_reg  (.CLK(clknet_leaf_151_clk_i_regs),
    .RESET_B(net1583),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_019_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_392_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[2]_reg  (.CLK(clknet_leaf_148_clk_i_regs),
    .RESET_B(net1562),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_020_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_391_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[30]_reg  (.CLK(clknet_leaf_152_clk_i_regs),
    .RESET_B(net1583),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_021_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_390_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[31]_reg  (.CLK(clknet_leaf_150_clk_i_regs),
    .RESET_B(net1582),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_022_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_389_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[3]_reg  (.CLK(clknet_leaf_148_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_023_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_388_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[4]_reg  (.CLK(clknet_leaf_148_clk_i_regs),
    .RESET_B(net1560),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_024_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_387_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[5]_reg  (.CLK(clknet_leaf_148_clk_i_regs),
    .RESET_B(net1562),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_025_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_386_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[6]_reg  (.CLK(clknet_leaf_147_clk_i_regs),
    .RESET_B(net1560),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_026_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_385_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[7]_reg  (.RESET_B(net1644),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_027_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [7]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_384_ ),
    .CLK(clknet_leaf_156_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[8]_reg  (.CLK(clknet_leaf_146_clk_i_regs),
    .RESET_B(net1644),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_028_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_383_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q[9]_reg  (.CLK(clknet_leaf_146_clk_i_regs),
    .RESET_B(net1644),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_029_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_414_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fetch_addr_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout473 (.A(\i_ibex/cs_registers_i/_0070_ ),
    .X(net473),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout472 (.A(\i_ibex/ex_block_i/alu_adder_result_ext [1]),
    .X(net472),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_530_  (.A(net703),
    .B_N(net1699),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_132_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_531_  (.A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy [0]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [1]),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_132_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_133_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_532_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_134_ ),
    .A(net698),
    .VSS(VSS));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_534_  (.B(net1471),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry_$_AND__Y_1_A ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_535_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_134_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_136_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_536_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_138_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_537_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .B(net1471),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_139_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_538_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .A2(net1471),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_140_ ),
    .B1(net698));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_539_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_141_ ),
    .A(instr_rdata_i[17]),
    .B(instr_rdata_i[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_540_  (.A(instr_err_i),
    .B(net1471),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_541_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_143_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [17]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_542_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .B_N(net1471),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_144_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(net472),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_544_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_146_ ),
    .A(net1478),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_545_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_144_ ),
    .C1(net1443),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_143_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_141_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_147_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_142_ ));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_546_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_139_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_140_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_147_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_547_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_149_ ),
    .A(instr_rdata_i[1]),
    .B(instr_rdata_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_548_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [1]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [0]),
    .A(net1470),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_549_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_150_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_151_ ),
    .VSS(VSS),
    .A1(net1470),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_149_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_550_  (.A0(net1699),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .S(net1470),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_152_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(net472),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_552_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_154_ ),
    .B(net1443),
    .A_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_152_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_553_  (.B1(\i_ibex/id_in_ready ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_155_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_151_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_154_ ));
 sg13g2_or2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_554_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_155_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(net472),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_556_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_137_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_138_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(net472),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout466 (.A(\i_ibex/cs_registers_i/_0037_ ),
    .X(net466),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_559_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_133_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout465 (.A(\i_ibex/cs_registers_i/_0037_ ),
    .X(net465),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout464 (.A(\i_ibex/cs_registers_i/_0037_ ),
    .X(net464),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_562_  (.A0(net1699),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [2]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_563_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ),
    .B(net1517),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_164_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_564_  (.B(net703),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry_$_AND__Y_A ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout463 (.A(\i_ibex/cs_registers_i/_0046_ ),
    .X(net463),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_566_  (.A(net1479),
    .B_N(net1439),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_567_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_164_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_167_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_568_  (.A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_136_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_168_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout462 (.A(\i_ibex/cs_registers_i/_0046_ ),
    .X(net462),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(\i_ibex/cs_registers_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_571_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_163_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [1]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(\i_ibex/cs_registers_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_573_  (.A0(net1699),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [2]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_574_  (.B(\i_ibex/pc_if [4]),
    .C(\i_ibex/pc_if [2]),
    .A(\i_ibex/pc_if [3]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_173_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_575_  (.B(\i_ibex/pc_if [5]),
    .C(\i_ibex/pc_if [6]),
    .A(\i_ibex/pc_if [7]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_174_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/pc_if [8]));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_576_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_175_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_174_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_173_ ));
 sg13g2_nor3_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_577_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ),
    .B(net1517),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_175_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(\i_ibex/cs_registers_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_579_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_178_ ),
    .A(\i_ibex/pc_if [9]),
    .B(net840),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_580_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_179_ ),
    .A(\i_ibex/pc_if [10]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(\i_ibex/cs_registers_i/_0079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_582_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_181_ ),
    .A(net1122),
    .VSS(VSS));
 sg13g2_buf_2 fanout457 (.A(\i_ibex/cs_registers_i/_0087_ ),
    .X(net457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(\i_ibex/cs_registers_i/_0087_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_585_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [10]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_179_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_586_  (.A(\i_ibex/pc_if [9]),
    .B(\i_ibex/pc_if [10]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_587_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_185_ ),
    .A(net840),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_184_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_588_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_186_ ),
    .A(\i_ibex/pc_if [11]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_589_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [11]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_186_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_590_  (.B(net1077),
    .C(net840),
    .A(\i_ibex/pc_if [11]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_187_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_184_ ));
 sg13g2_buf_2 fanout455 (.A(\i_ibex/cs_registers_i/_0104_ ),
    .X(net455),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_592_  (.A0(\i_ibex/pc_if [12]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [12]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_593_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_005_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_187_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_594_  (.B(\i_ibex/pc_if [10]),
    .C(\i_ibex/pc_if [12]),
    .A(\i_ibex/pc_if [9]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_190_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/pc_if [11]));
 sg13g2_nor3_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_595_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_175_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_190_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_596_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .A(\i_ibex/pc_if [13]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_192_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_597_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [13]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_192_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_598_  (.B(\i_ibex/pc_if [13]),
    .A(\i_ibex/pc_if [14]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_599_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_194_ ),
    .B(net1115),
    .A_N(\i_ibex/if_stage_i/fetch_addr_n [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_600_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_194_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_195_ ),
    .VSS(VSS),
    .A1(net1128),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_193_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_601_  (.A0(\i_ibex/pc_if [14]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [14]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_602_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_196_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_197_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_603_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_195_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_007_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_197_ ));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_604_  (.A(net1115),
    .B_N(\i_ibex/pc_if [15]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_198_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_605_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1115),
    .A2(\i_ibex/if_stage_i/fetch_addr_n [15]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_199_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_198_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_606_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_200_ ),
    .A(\i_ibex/pc_if [14]),
    .B(\i_ibex/pc_if [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_607_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_201_ ),
    .A(\i_ibex/pc_if [15]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_608_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [15]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_201_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_609_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_203_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_610_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_203_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_008_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_199_ ));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_611_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_204_ ),
    .A(\i_ibex/pc_if [16]),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_612_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_205_ ),
    .A(net1115),
    .B(\i_ibex/if_stage_i/fetch_addr_n [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_613_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_205_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_206_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_204_ ),
    .A2(net1122));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_614_  (.B(\i_ibex/pc_if [14]),
    .C(\i_ibex/pc_if [13]),
    .A(\i_ibex/pc_if [15]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_615_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_208_ ),
    .A(\i_ibex/pc_if [16]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_616_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [16]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_208_ ),
    .S(net1078),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_209_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_617_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_206_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_209_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_191_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_618_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_204_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_190_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_207_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_210_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_619_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_211_ ),
    .A(net839),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_210_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_620_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_212_ ),
    .A(\i_ibex/pc_if [17]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_621_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [17]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_212_ ),
    .S(net1075),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_622_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_213_ ),
    .A(\i_ibex/pc_if [17]),
    .B(net839),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_210_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_623_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_213_ ),
    .A(\i_ibex/pc_if [18]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_214_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_624_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [18]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_214_ ),
    .S(net1075),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_625_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_215_ ),
    .A(\i_ibex/pc_if [18]),
    .B(\i_ibex/pc_if [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_626_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_204_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_190_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_207_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_215_ ));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_627_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_217_ ),
    .A(net839),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_628_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_218_ ),
    .A(\i_ibex/pc_if [19]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_217_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_629_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [19]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_218_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_630_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_219_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_154_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_151_ ));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_632_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_221_ ),
    .B(net1470),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_633_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_222_ ),
    .A(\i_ibex/id_in_ready ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_221_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_634_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_223_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_143_ ),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_144_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_142_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_635_  (.B1(net1477),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_224_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_223_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_222_ ));
 sg13g2_o21ai_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_636_  (.B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_224_ ),
    .VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ),
    .VSS(VSS),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_219_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_222_ ));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(net455),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_638_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [1]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ),
    .S(net1078),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_639_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_227_ ),
    .A(\i_ibex/pc_if [19]),
    .B(net1074),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_640_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_228_ ),
    .A(net839),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_227_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_641_  (.A0(\i_ibex/pc_if [20]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [20]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_229_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_642_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_014_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_228_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_229_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_643_  (.A(\i_ibex/pc_if [20]),
    .B(\i_ibex/pc_if [19]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_230_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_644_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_230_ ),
    .A(net838),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_645_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_232_ ),
    .A(\i_ibex/pc_if [21]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_231_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_646_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [21]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_232_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_647_  (.B(net838),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .A(\i_ibex/pc_if [21]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_230_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_648_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_234_ ),
    .A(\i_ibex/pc_if [22]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_233_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_649_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [22]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_234_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_650_  (.A(\i_ibex/pc_if [22]),
    .B(\i_ibex/pc_if [21]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_235_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_651_  (.B(net838),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_227_ ),
    .A(\i_ibex/pc_if [20]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_236_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_235_ ));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_652_  (.A0(\i_ibex/pc_if [23]),
    .A1(\i_ibex/if_stage_i/fetch_addr_n [23]),
    .S(net1140),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_653_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_017_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_236_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_237_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_654_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_238_ ),
    .A(\i_ibex/pc_if [23]),
    .B(\i_ibex/pc_if [22]),
    .C(\i_ibex/pc_if [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_655_  (.A(net838),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_230_ ),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_238_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_239_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_656_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_239_ ),
    .A(\i_ibex/pc_if [24]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_240_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_657_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [24]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_240_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_658_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_241_ ),
    .A(\i_ibex/pc_if [24]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_230_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_238_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_659_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_241_ ),
    .A(net838),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_660_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_243_ ),
    .A(\i_ibex/pc_if [25]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_661_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [25]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_243_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_662_  (.X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_244_ ),
    .A(\i_ibex/pc_if [25]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_241_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_663_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_245_ ),
    .A(net838),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_664_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_246_ ),
    .A(\i_ibex/pc_if [26]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_245_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_665_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [26]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_246_ ),
    .S(net1075),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_666_  (.B(net838),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_244_ ),
    .A(\i_ibex/pc_if [26]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_667_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_248_ ),
    .A(\i_ibex/pc_if [27]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_247_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_668_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [27]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_248_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_669_  (.B(\i_ibex/pc_if [26]),
    .C(net838),
    .A(\i_ibex/pc_if [27]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_249_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_244_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_670_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_250_ ),
    .A(\i_ibex/pc_if [28]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_249_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_671_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [28]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_250_ ),
    .S(net1075),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_672_  (.B(\i_ibex/pc_if [26]),
    .C(\i_ibex/pc_if [28]),
    .A(\i_ibex/pc_if [27]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_251_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_673_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_174_ ),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_251_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_252_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_674_  (.B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_216_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_241_ ),
    .A(\i_ibex/pc_if [25]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_253_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_252_ ));
 sg13g2_nor4_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_675_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ),
    .B(net1517),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_173_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_253_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_676_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_255_ ),
    .A(\i_ibex/pc_if [29]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_677_  (.A(net1076),
    .B(\i_ibex/if_stage_i/fetch_addr_n [29]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_256_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_678_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1076),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_255_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_023_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_256_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_679_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_257_ ),
    .A(\i_ibex/pc_if [2]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_680_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [2]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_257_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_681_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_258_ ),
    .A(\i_ibex/pc_if [29]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_254_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_682_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_259_ ),
    .A(\i_ibex/pc_if [30]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_258_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_683_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [30]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_259_ ),
    .S(net1074),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_684_  (.B(\i_ibex/pc_if [30]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_254_ ),
    .A(\i_ibex/pc_if [29]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_685_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_261_ ),
    .A(\i_ibex/pc_if [31]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_260_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_686_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [31]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_261_ ),
    .S(net1076),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_687_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_262_ ),
    .A(\i_ibex/pc_if [2]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_164_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_688_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_263_ ),
    .A(\i_ibex/pc_if [3]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_262_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_689_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [3]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_263_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_690_  (.B(\i_ibex/pc_if [2]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_164_ ),
    .A(\i_ibex/pc_if [3]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_691_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_265_ ),
    .A(\i_ibex/pc_if [4]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_264_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_692_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [4]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_265_ ),
    .S(net1077),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_693_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ),
    .B(net1517),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_173_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_694_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_267_ ),
    .A(\i_ibex/pc_if [5]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_695_  (.A(net1079),
    .B(\i_ibex/if_stage_i/fetch_addr_n [5]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_268_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_696_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net1079),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_267_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_029_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_268_ ));
 sg13g2_nand2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_697_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_269_ ),
    .A(\i_ibex/pc_if [5]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_266_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_698_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_270_ ),
    .A(\i_ibex/pc_if [6]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_269_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_699_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [6]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_270_ ),
    .S(net1079),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_700_  (.B(\i_ibex/pc_if [6]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_266_ ),
    .A(\i_ibex/pc_if [5]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_271_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_701_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_272_ ),
    .A(\i_ibex/pc_if [7]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_271_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_702_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [7]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_272_ ),
    .S(net1079),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_703_  (.B(\i_ibex/pc_if [5]),
    .C(\i_ibex/pc_if [6]),
    .A(\i_ibex/pc_if [7]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_273_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_266_ ));
 sg13g2_xnor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_704_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_274_ ),
    .A(\i_ibex/pc_if [8]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_273_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_705_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [8]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_274_ ),
    .S(net1079),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_706_  (.B(net840),
    .A(\i_ibex/pc_if [9]),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_275_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_707_  (.A0(\i_ibex/if_stage_i/fetch_addr_n [9]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_275_ ),
    .S(net1076),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout452 (.A(\i_ibex/ex_block_i/alu_i/_0677_ ),
    .X(net452),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_709_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .B(net1471),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_277_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_710_  (.A(instr_err_i),
    .B(net703),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_277_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_278_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_711_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [1]),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_134_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_279_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_712_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_280_ ),
    .B(net698),
    .A(net1470));
 sg13g2_a221oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_713_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .C1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_223_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_280_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_134_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_281_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry [0]));
 sg13g2_nor4_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_714_  (.A(net1443),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_278_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_279_ ),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_281_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_282_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_715_  (.A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_152_ ),
    .A1(net1443),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_282_ ),
    .X(\i_ibex/if_stage_i/fetch_err ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_716_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_283_ ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_plus2_$_AND__Y_B ),
    .VSS(VSS));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(\i_ibex/cs_registers_i/_0129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_718_  (.Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_285_ ),
    .B1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_132_ ),
    .B2(net1471),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy [0]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_719_  (.A(net1443),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_283_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_285_ ),
    .Y(\i_ibex/if_stage_i/fetch_err_plus2 ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(\i_ibex/cs_registers_i/_0129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_721_  (.A0(net1681),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [47]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_287_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout449 (.A(\i_ibex/cs_registers_i/_0136_ ),
    .X(net449),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_723_  (.A0(instr_rdata_i[31]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [31]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_289_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_724_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_287_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_289_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_725_  (.A0(net1684),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [46]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_290_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_726_  (.A0(net1703),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [30]),
    .S(net1472),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_291_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_727_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_290_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_291_ ),
    .S(net1443),
    .X(\i_ibex/if_stage_i/fetch_rdata [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(\i_ibex/cs_registers_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_729_  (.A0(net1735),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [37]),
    .S(net702),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_293_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_730_  (.A0(instr_rdata_i[21]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [21]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_294_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_731_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_293_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_294_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_732_  (.A0(net1679),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [36]),
    .S(net702),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_295_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_733_  (.A0(net1697),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [20]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_734_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_295_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_296_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_735_  (.A0(net1675),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [35]),
    .S(net702),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_297_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_736_  (.A0(instr_rdata_i[19]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [19]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_298_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_737_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_297_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_298_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_738_  (.A0(net1719),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [34]),
    .S(net702),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_299_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_739_  (.A0(instr_rdata_i[18]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [18]),
    .S(net1475),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_300_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_740_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_299_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_300_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_741_  (.A0(net1691),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [33]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_301_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_742_  (.A0(instr_rdata_i[17]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [17]),
    .S(net1472),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_743_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_301_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_302_ ),
    .S(net1444),
    .X(\i_ibex/if_stage_i/fetch_rdata [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_744_  (.A0(net1698),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [32]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_303_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_745_  (.A0(instr_rdata_i[16]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [16]),
    .S(net1472),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_304_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_746_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_303_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_304_ ),
    .S(net1443),
    .X(\i_ibex/if_stage_i/fetch_rdata [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_747_  (.A0(instr_rdata_i[15]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [15]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(\i_ibex/cs_registers_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_749_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_289_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_305_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_750_  (.A0(instr_rdata_i[14]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [14]),
    .S(net1470),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_307_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_751_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_291_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_307_ ),
    .S(net1444),
    .X(\i_ibex/if_stage_i/fetch_rdata [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(\i_ibex/cs_registers_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_753_  (.A0(instr_rdata_i[29]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [29]),
    .S(net1475),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_309_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_754_  (.A0(instr_rdata_i[13]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [13]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_755_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_309_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_310_ ),
    .S(net1447),
    .X(\i_ibex/if_stage_i/fetch_rdata [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_756_  (.A0(net1674),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [28]),
    .S(net1475),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_311_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_757_  (.A0(instr_rdata_i[12]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [12]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_312_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_758_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_311_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_312_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_759_  (.A0(net1708),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [45]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_760_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_309_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_313_ ),
    .S(net1478),
    .X(\i_ibex/if_stage_i/fetch_rdata [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_761_  (.A0(instr_rdata_i[27]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [27]),
    .S(net1475),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_314_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_762_  (.A0(instr_rdata_i[11]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [11]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_763_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_314_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_315_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_764_  (.A0(instr_rdata_i[26]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [26]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_316_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_765_  (.A0(net1710),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [10]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_317_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_766_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_316_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_317_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_767_  (.A0(net1683),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [25]),
    .S(net1471),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_318_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_768_  (.A0(net1724),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [9]),
    .S(net1470),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_319_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_769_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_318_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_319_ ),
    .S(net1444),
    .X(\i_ibex/if_stage_i/fetch_rdata [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_770_  (.A0(net1693),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [24]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_320_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_771_  (.A0(net1688),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [8]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_321_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_772_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_320_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_321_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_773_  (.A0(instr_rdata_i[23]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [23]),
    .S(net1475),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_322_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_774_  (.A0(net1696),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [7]),
    .S(net1476),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_775_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_322_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_323_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_776_  (.A0(net1680),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [22]),
    .S(net1474),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_324_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_777_  (.A0(net1689),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [6]),
    .S(net1476),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_325_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_778_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_324_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_325_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_779_  (.A0(net1735),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [5]),
    .S(net1476),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_326_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_780_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_294_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_326_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_781_  (.A0(net1679),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [4]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_327_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_782_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_296_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_327_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_783_  (.A0(net1675),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [3]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_328_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_784_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_298_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_328_ ),
    .S(net1446),
    .X(\i_ibex/if_stage_i/fetch_rdata [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_785_  (.A0(net1719),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [2]),
    .S(net1473),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_786_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_300_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_329_ ),
    .S(net1445),
    .X(\i_ibex/if_stage_i/fetch_rdata [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_787_  (.A0(net1702),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [44]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_330_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_788_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_311_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_330_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_789_  (.A0(instr_rdata_i[1]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [1]),
    .S(net1472),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_331_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_790_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_302_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_331_ ),
    .S(net1444),
    .X(\i_ibex/if_stage_i/fetch_rdata [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_791_  (.A0(instr_rdata_i[0]),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [0]),
    .S(net1472),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_332_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_792_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_304_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_332_ ),
    .S(net1443),
    .X(\i_ibex/if_stage_i/fetch_rdata [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_793_  (.A0(net1687),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [43]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_333_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_794_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_314_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_333_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_795_  (.A0(net1710),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [42]),
    .S(net701),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_334_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_796_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_316_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_334_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_797_  (.A0(net1724),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [41]),
    .S(net698),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_335_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_798_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_318_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_335_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_799_  (.A0(net1688),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [40]),
    .S(net698),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_800_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_320_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_336_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_801_  (.A0(net1696),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [39]),
    .S(net698),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_337_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_802_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_322_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_337_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_803_  (.A0(net1689),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [38]),
    .S(net698),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_338_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_804_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_324_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_338_ ),
    .S(net1477),
    .X(\i_ibex/if_stage_i/fetch_rdata [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_805_  (.VDD(VDD),
    .Y(\i_ibex/if_stage_i/fetch_valid ),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_806_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_303_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [0]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_807_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_334_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [10]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_808_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_333_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [11]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_809_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_330_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [12]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_810_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_313_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [13]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_811_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_290_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [14]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_812_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_287_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [15]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_040_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_813_  (.A0(net1709),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [48]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_339_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_814_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_339_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [16]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_041_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_815_  (.A0(net1676),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [49]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_340_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_816_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_340_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [17]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_817_  (.A0(net1678),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [50]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_341_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(\i_ibex/cs_registers_i/_0161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_819_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_341_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [18]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_820_  (.A0(net1690),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [51]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_343_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_821_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_343_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [19]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_822_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_301_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [1]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_823_  (.A0(net1697),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [52]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_344_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_824_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_344_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [20]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_825_  (.A0(net1682),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [53]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_345_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_826_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_345_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [21]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_827_  (.A0(net1680),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [54]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_346_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_828_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_346_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [22]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_829_  (.A0(net1686),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [55]),
    .S(net699),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_347_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_830_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_347_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [23]),
    .S(net816),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_831_  (.A0(net1693),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [56]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_348_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_832_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_348_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [24]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_833_  (.A0(net1683),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [57]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_349_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_834_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_349_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [25]),
    .S(net816),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_835_  (.A0(net1692),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [58]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_350_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_836_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_350_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [26]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_837_  (.A0(net1700),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [59]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_351_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout444 (.A(\i_ibex/ex_block_i/alu_i/_0083_ ),
    .X(net444),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_839_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_351_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [27]),
    .S(net816),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_840_  (.A0(net1674),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [60]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_353_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_841_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_353_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [28]),
    .S(net818),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_842_  (.A0(net1685),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [61]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_354_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_843_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_354_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [29]),
    .S(net819),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_844_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_299_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [2]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_845_  (.A0(net1703),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [62]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_355_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_846_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_355_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [30]),
    .S(net816),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_847_  (.A0(net1701),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [63]),
    .S(net700),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_356_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_848_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_356_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [31]),
    .S(net819),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_058_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_849_  (.A0(net1698),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [64]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_357_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_850_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_357_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [32]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_851_  (.A0(net1691),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [65]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_358_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_852_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_358_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [33]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_060_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_853_  (.A0(net1719),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [66]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_359_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_854_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_359_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [34]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_855_  (.A0(net1675),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [67]),
    .S(net1483),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_360_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_856_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_360_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [35]),
    .S(net814),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_857_  (.A0(net1679),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [68]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_361_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_858_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_361_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [36]),
    .S(net814),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_859_  (.A0(net1735),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [69]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_362_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_860_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_362_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [37]),
    .S(net814),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_064_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_861_  (.A0(net1689),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [70]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_363_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_862_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_363_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [38]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_863_  (.A0(net1696),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [71]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_364_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_864_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_364_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [39]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_066_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_865_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_297_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [3]),
    .S(net819),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_067_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_866_  (.A0(net1688),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [72]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_365_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_867_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_365_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [40]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_068_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout443 (.A(net444),
    .X(net443),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_869_  (.A0(net1724),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [73]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_367_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout442 (.A(net444),
    .X(net442),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_871_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_367_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [41]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_872_  (.A0(net1710),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [74]),
    .S(net1483),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_369_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_873_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_369_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [42]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_070_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_874_  (.A0(net1687),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [75]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_370_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_875_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_370_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [43]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_071_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_876_  (.A0(net1702),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [76]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_371_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_877_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_371_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [44]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_072_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_878_  (.A0(net1708),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [77]),
    .S(net1481),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_372_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_879_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_372_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [45]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_073_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_880_  (.A0(net1684),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [78]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_373_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_881_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_373_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [46]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_074_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_882_  (.A0(net1681),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [79]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_374_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_883_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_374_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [47]),
    .S(net812),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_075_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_884_  (.A0(net1709),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [80]),
    .S(net1480),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_375_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_885_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_375_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [48]),
    .S(net811),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_076_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_886_  (.A0(net1676),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [81]),
    .S(net1480),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_376_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_887_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_376_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [49]),
    .S(net811),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_077_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_888_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_295_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [4]),
    .S(net819),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_889_  (.A0(net1678),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [82]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_377_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_890_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_377_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [50]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_079_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout441 (.A(net444),
    .X(net441),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_892_  (.A0(net1690),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [83]),
    .S(net1483),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_379_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout440 (.A(\i_ibex/ex_block_i/alu_i/_0083_ ),
    .X(net440),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_894_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_379_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [51]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_895_  (.A0(net1697),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [84]),
    .S(net1483),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_381_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_896_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_381_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [52]),
    .S(net814),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_081_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_897_  (.A0(net1682),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [85]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_382_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_898_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_382_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [53]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_899_  (.A0(net1680),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [86]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_383_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_900_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_383_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [54]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_083_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_901_  (.A0(net1686),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [87]),
    .S(net1480),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_384_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_902_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_384_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [55]),
    .S(net811),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_084_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_903_  (.A0(net1693),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [88]),
    .S(net1483),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_385_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_904_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_385_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [56]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_085_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_905_  (.A0(net1683),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [89]),
    .S(net1480),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_386_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_906_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_386_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [57]),
    .S(net811),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_086_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_907_  (.A0(net1692),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [90]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_387_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_908_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_387_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [58]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_087_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_909_  (.A0(net1700),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [91]),
    .S(net1480),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_388_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_910_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_388_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [59]),
    .S(net811),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_911_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_293_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [5]),
    .S(net819),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_089_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_912_  (.A0(net1674),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [92]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_389_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_913_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_389_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [60]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_090_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_914_  (.A0(net1685),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [93]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_915_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_390_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [61]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_091_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_916_  (.A0(net1703),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [94]),
    .S(net1479),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_391_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_917_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_391_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [62]),
    .S(net810),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_918_  (.A0(net1701),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [95]),
    .S(net1482),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_392_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_919_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_392_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [63]),
    .S(net813),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_920_  (.A0(net1698),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [64]),
    .S(net1439),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_094_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_921_  (.A0(net1691),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [65]),
    .S(net1439),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_095_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_922_  (.A0(net1719),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [66]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_096_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_923_  (.A0(net1675),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [67]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_924_  (.A0(net1679),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [68]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_098_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_925_  (.A0(net1735),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [69]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_099_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_926_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_338_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [6]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_100_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_927_  (.A0(net1689),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [70]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_101_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_928_  (.A0(net1696),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [71]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_102_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_929_  (.A0(net1688),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [72]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout439 (.A(net440),
    .X(net439),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_931_  (.A0(net1724),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [73]),
    .S(net1439),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_104_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_932_  (.A0(net1710),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [74]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_933_  (.A0(net1687),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [75]),
    .S(net1439),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_106_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_934_  (.A0(net1702),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [76]),
    .S(net1439),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_107_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_935_  (.A0(net1708),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [77]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_108_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_936_  (.A0(net1684),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [78]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_109_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_937_  (.A0(net1681),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [79]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_938_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_337_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [7]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_111_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_939_  (.A0(net1709),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [80]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_940_  (.A0(net1676),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [81]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_941_  (.A0(net1678),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [82]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_114_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(net440),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_943_  (.A0(net1690),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [83]),
    .S(net1442),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_944_  (.A0(net1697),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [84]),
    .S(net1442),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_116_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_945_  (.A0(net1682),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [85]),
    .S(net1442),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_117_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_946_  (.A0(net1680),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [86]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_118_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_947_  (.A0(net1686),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [87]),
    .S(net1439),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_119_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_948_  (.A0(net1693),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [88]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_120_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_949_  (.A0(net1683),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [89]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_121_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_950_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_336_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [8]),
    .S(net817),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_951_  (.A0(net1692),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [90]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_123_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_952_  (.A0(net1700),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [91]),
    .S(net1442),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_124_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_953_  (.A0(net1674),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [92]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_954_  (.A0(net1685),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [93]),
    .S(net1441),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_126_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_955_  (.A0(net1703),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [94]),
    .S(net1438),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_127_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_956_  (.A0(net1701),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [95]),
    .S(net1440),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_957_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_335_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [9]),
    .S(net815),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_958_  (.A(net1126),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_164_ ),
    .C(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_167_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_959_  (.VSS(VSS),
    .VDD(VDD),
    .B1(net1126),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_395_ ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_137_ ));
 sg13g2_nor2b_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_960_  (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_168_ ),
    .B_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_395_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_961_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_valid ),
    .A2(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry [0]),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_396_ ),
    .B1(net1470));
 sg13g2_mux2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_962_  (.A0(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_137_ ),
    .A1(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_396_ ),
    .S(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_156_ ),
    .X(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_397_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_963_  (.A(net1126),
    .B(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_397_ ),
    .Y(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(net1051),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/busy_o[0]_reg  (.CLK(clknet_leaf_112_clk_i_regs),
    .RESET_B(net1663),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d [1]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry_$_AND__Y_1_A ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/busy_o[1]_reg  (.CLK(clknet_leaf_112_clk_i_regs),
    .RESET_B(net1663),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d [2]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry_$_AND__Y_A ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_000_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [0]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_plus2_$_AND__Y_B ),
    .CLK(clknet_leaf_113_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q[1]_reg  (.CLK(clknet_leaf_113_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_001_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_525_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q[2]_reg  (.CLK(clknet_leaf_113_clk_i_regs),
    .RESET_B(net1663),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_002_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_524_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/err_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[10]_reg  (.RESET_B(net1584),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_003_ ),
    .Q(\i_ibex/pc_if [10]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_523_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[11]_reg  (.RESET_B(net1583),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_004_ ),
    .Q(\i_ibex/pc_if [11]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_522_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[12]_reg  (.RESET_B(net1582),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_005_ ),
    .Q(\i_ibex/pc_if [12]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_521_ ),
    .CLK(clknet_leaf_140_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[13]_reg  (.RESET_B(net1584),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_006_ ),
    .Q(\i_ibex/pc_if [13]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_520_ ),
    .CLK(clknet_leaf_142_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[14]_reg  (.RESET_B(net1582),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_007_ ),
    .Q(\i_ibex/pc_if [14]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_519_ ),
    .CLK(clknet_leaf_149_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[15]_reg  (.RESET_B(net1582),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_008_ ),
    .Q(\i_ibex/pc_if [15]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_518_ ),
    .CLK(clknet_leaf_142_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[16]_reg  (.RESET_B(net1582),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_009_ ),
    .Q(\i_ibex/pc_if [16]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_517_ ),
    .CLK(clknet_leaf_142_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[17]_reg  (.RESET_B(net1625),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_010_ ),
    .Q(\i_ibex/pc_if [17]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_516_ ),
    .CLK(clknet_leaf_150_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[18]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_011_ ),
    .Q(\i_ibex/pc_if [18]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_515_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[19]_reg  (.RESET_B(net1646),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_012_ ),
    .Q(\i_ibex/pc_if [19]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_514_ ),
    .CLK(clknet_leaf_151_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[1]_reg  (.CLK(clknet_leaf_84_clk_i_regs),
    .RESET_B(net1610),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_013_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_513_ ),
    .Q(\i_ibex/pc_if [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[20]_reg  (.RESET_B(net1645),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_014_ ),
    .Q(\i_ibex/pc_if [20]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_512_ ),
    .CLK(clknet_leaf_151_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[21]_reg  (.RESET_B(net1645),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_015_ ),
    .Q(\i_ibex/pc_if [21]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_511_ ),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[22]_reg  (.RESET_B(net1645),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_016_ ),
    .Q(\i_ibex/pc_if [22]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_510_ ),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[23]_reg  (.RESET_B(net1646),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_017_ ),
    .Q(\i_ibex/pc_if [23]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_509_ ),
    .CLK(clknet_leaf_151_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[24]_reg  (.RESET_B(net1646),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_018_ ),
    .Q(\i_ibex/pc_if [24]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_508_ ),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[25]_reg  (.RESET_B(net1625),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_019_ ),
    .Q(\i_ibex/pc_if [25]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_507_ ),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[26]_reg  (.RESET_B(net1625),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_020_ ),
    .Q(\i_ibex/pc_if [26]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_506_ ),
    .CLK(clknet_leaf_151_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[27]_reg  (.RESET_B(net1625),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_021_ ),
    .Q(\i_ibex/pc_if [27]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_505_ ),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[28]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_022_ ),
    .Q(\i_ibex/pc_if [28]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_504_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[29]_reg  (.RESET_B(net1627),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_023_ ),
    .Q(\i_ibex/pc_if [29]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_503_ ),
    .CLK(clknet_leaf_139_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[2]_reg  (.RESET_B(net1610),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_024_ ),
    .Q(\i_ibex/pc_if [2]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_502_ ),
    .CLK(clknet_leaf_82_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[30]_reg  (.RESET_B(net1625),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_025_ ),
    .Q(\i_ibex/pc_if [30]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_501_ ),
    .CLK(clknet_leaf_140_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[31]_reg  (.RESET_B(net1626),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_026_ ),
    .Q(\i_ibex/pc_if [31]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_500_ ),
    .CLK(clknet_leaf_139_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[3]_reg  (.RESET_B(net1610),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_027_ ),
    .Q(\i_ibex/pc_if [3]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_499_ ),
    .CLK(clknet_leaf_82_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[4]_reg  (.RESET_B(net1610),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_028_ ),
    .Q(\i_ibex/pc_if [4]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_498_ ),
    .CLK(clknet_leaf_82_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[5]_reg  (.RESET_B(net1606),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_029_ ),
    .Q(\i_ibex/pc_if [5]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_497_ ),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[6]_reg  (.RESET_B(net1567),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_030_ ),
    .Q(\i_ibex/pc_if [6]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_496_ ),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[7]_reg  (.RESET_B(net1567),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_031_ ),
    .Q(\i_ibex/pc_if [7]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_495_ ),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[8]_reg  (.RESET_B(net1567),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_032_ ),
    .Q(\i_ibex/pc_if [8]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_494_ ),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/out_addr_o[9]_reg  (.RESET_B(net1582),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_033_ ),
    .Q(\i_ibex/pc_if [9]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_493_ ),
    .CLK(clknet_leaf_141_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[0]_reg  (.CLK(clknet_leaf_113_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_034_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_492_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[10]_reg  (.CLK(clknet_leaf_125_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_035_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_491_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[11]_reg  (.CLK(clknet_leaf_116_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_036_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_490_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[12]_reg  (.CLK(clknet_leaf_120_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_037_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_489_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[13]_reg  (.CLK(clknet_5_20__leaf_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_038_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_488_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[14]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_039_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_487_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[15]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_040_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_486_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[16]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_041_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_485_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[17]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_042_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_484_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[18]_reg  (.CLK(clknet_leaf_118_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_043_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_483_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[19]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_044_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_482_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[1]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_045_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_481_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[20]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_046_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_480_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[21]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_047_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_479_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[22]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_048_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_478_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[23]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_049_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_477_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[24]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_050_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_476_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[25]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(net1663),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_051_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_475_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[26]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_052_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_474_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[27]_reg  (.CLK(clknet_leaf_116_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_053_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_473_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[28]_reg  (.CLK(clknet_leaf_118_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_054_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_472_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[29]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_055_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_471_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[2]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_056_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_470_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[30]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_057_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_469_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[31]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_058_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_468_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[32]_reg  (.CLK(clknet_leaf_113_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_059_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_467_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [32]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[33]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_060_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_466_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [33]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[34]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_061_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_465_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [34]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[35]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_062_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_464_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [35]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[36]_reg  (.CLK(clknet_leaf_120_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_063_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_463_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [36]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[37]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_064_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_462_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [37]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[38]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_065_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_461_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [38]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[39]_reg  (.CLK(clknet_leaf_131_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_066_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_460_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [39]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[3]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_067_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_459_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[40]_reg  (.CLK(clknet_leaf_131_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_068_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_458_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [40]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[41]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_069_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_457_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [41]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[42]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_070_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_456_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [42]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[43]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_071_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_455_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [43]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[44]_reg  (.CLK(clknet_leaf_120_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_072_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_454_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [44]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[45]_reg  (.CLK(clknet_leaf_131_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_073_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_453_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [45]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[46]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_074_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_452_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [46]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[47]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_075_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_451_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [47]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[48]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_076_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_450_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [48]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[49]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_077_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_449_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [49]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[4]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_078_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_448_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[50]_reg  (.CLK(clknet_leaf_118_clk_i_regs),
    .RESET_B(net1662),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_079_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_447_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [50]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[51]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_080_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_446_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [51]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[52]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_081_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_445_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [52]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[53]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_082_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_444_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [53]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[54]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_083_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_443_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [54]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[55]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_084_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_442_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [55]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[56]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_085_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_441_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [56]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[57]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1661),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_086_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_440_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [57]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[58]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_087_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_439_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [58]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[59]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1661),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_088_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_438_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [59]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[5]_reg  (.CLK(clknet_leaf_126_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_089_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_437_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[60]_reg  (.CLK(clknet_leaf_118_clk_i_regs),
    .RESET_B(net1662),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_090_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_436_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [60]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[61]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_091_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_435_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [61]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[62]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(net1663),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_092_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_434_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [62]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[63]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_093_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_433_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [63]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[64]_reg  (.CLK(clknet_leaf_113_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_094_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_432_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [64]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[65]_reg  (.CLK(clknet_leaf_113_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_095_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_431_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [65]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[66]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_096_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_430_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [66]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[67]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_097_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_429_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [67]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[68]_reg  (.CLK(clknet_leaf_120_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_098_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_428_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [68]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[69]_reg  (.CLK(clknet_leaf_126_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_099_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_427_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [69]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[6]_reg  (.CLK(clknet_leaf_125_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_100_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_426_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[70]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_101_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_425_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [70]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[71]_reg  (.CLK(clknet_leaf_131_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_102_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_424_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [71]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[72]_reg  (.CLK(clknet_leaf_131_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_103_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_423_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [72]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[73]_reg  (.CLK(clknet_leaf_111_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_104_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_422_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [73]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[74]_reg  (.CLK(clknet_leaf_125_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_105_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_421_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [74]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[75]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_106_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_420_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [75]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[76]_reg  (.CLK(clknet_leaf_116_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_107_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_419_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [76]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[77]_reg  (.CLK(clknet_leaf_131_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_108_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_418_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [77]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[78]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_109_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_417_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [78]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[79]_reg  (.CLK(clknet_leaf_120_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_110_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_416_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [79]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[7]_reg  (.CLK(clknet_leaf_125_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_111_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_415_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[80]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_112_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_414_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [80]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[81]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1660),
    .D(net1677),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_413_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [81]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[82]_reg  (.CLK(clknet_leaf_118_clk_i_regs),
    .RESET_B(net1662),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_114_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_412_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [82]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[83]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(net1663),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_115_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_411_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [83]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[84]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_116_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_410_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [84]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[85]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_117_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_409_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [85]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[86]_reg  (.CLK(clknet_leaf_122_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_118_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_408_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [86]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[87]_reg  (.CLK(clknet_leaf_117_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_119_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_407_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [87]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[88]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_120_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_406_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [88]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[89]_reg  (.CLK(clknet_leaf_115_clk_i_regs),
    .RESET_B(net1661),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_121_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_405_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [89]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[8]_reg  (.CLK(clknet_leaf_124_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_122_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_404_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[90]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_123_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_403_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [90]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[91]_reg  (.CLK(clknet_leaf_116_clk_i_regs),
    .RESET_B(net1661),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_124_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_402_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [91]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[92]_reg  (.CLK(clknet_leaf_119_clk_i_regs),
    .RESET_B(net1662),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_125_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_401_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [92]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[93]_reg  (.CLK(clknet_leaf_121_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_126_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_400_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [93]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[94]_reg  (.CLK(clknet_leaf_114_clk_i_regs),
    .RESET_B(net1660),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_127_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_399_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [94]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[95]_reg  (.CLK(clknet_leaf_123_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_128_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_398_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [95]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q[9]_reg  (.CLK(clknet_leaf_111_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_129_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_526_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/rdata_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_q[0]_reg  (.CLK(clknet_leaf_112_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_d [0]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/lowest_free_entry [0]),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q[0]_reg  (.CLK(clknet_leaf_142_clk_i_regs),
    .RESET_B(net1562),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_s [0]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_415_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q[1]_reg  (.CLK(clknet_leaf_143_clk_i_regs),
    .RESET_B(net1562),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_s [1]),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__Y_B ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/rdata_outstanding_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[10]_reg  (.CLK(clknet_leaf_146_clk_i_regs),
    .RESET_B(net1644),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_030_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_382_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[11]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_031_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_381_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[12]_reg  (.CLK(clknet_leaf_144_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_032_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_380_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[13]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1641),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_033_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_379_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[14]_reg  (.CLK(clknet_leaf_148_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_034_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_378_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[15]_reg  (.CLK(clknet_leaf_144_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_035_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_377_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[16]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1561),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_036_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_376_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[17]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1641),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_037_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_375_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[18]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_038_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_374_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[19]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_039_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_373_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[20]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_040_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_372_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[21]_reg  (.CLK(clknet_leaf_4_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_041_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_371_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[22]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_042_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_370_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[23]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1647),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_043_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_369_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[24]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_044_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_368_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[25]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1638),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_045_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_367_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[26]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1641),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_046_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_366_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[27]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_047_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_365_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[28]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1643),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_048_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_364_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[29]_reg  (.CLK(clknet_leaf_2_clk_i_regs),
    .RESET_B(net1640),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_049_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_363_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[2]_reg  (.CLK(clknet_leaf_143_clk_i_regs),
    .RESET_B(net1652),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_050_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_362_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[30]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1561),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_051_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_361_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[31]_reg  (.CLK(clknet_leaf_146_clk_i_regs),
    .RESET_B(net1644),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_052_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_360_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[3]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1641),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_053_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_359_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[4]_reg  (.CLK(clknet_leaf_144_clk_i_regs),
    .RESET_B(net1651),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_054_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_358_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[5]_reg  (.CLK(clknet_leaf_144_clk_i_regs),
    .RESET_B(net1652),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_055_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_357_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[6]_reg  (.CLK(clknet_leaf_155_clk_i_regs),
    .RESET_B(net1642),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_056_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_356_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[7]_reg  (.CLK(clknet_leaf_154_clk_i_regs),
    .RESET_B(net1641),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_057_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_355_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[8]_reg  (.CLK(clknet_leaf_156_clk_i_regs),
    .RESET_B(net1644),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_058_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_354_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q[9]_reg  (.CLK(clknet_leaf_146_clk_i_regs),
    .RESET_B(net1644),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/_059_ ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/_416_ ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/stored_addr_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/if_stage_i/prefetch_buffer_i/valid_req_q_reg  (.RESET_B(net1651),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/if_stage_i/prefetch_buffer_i/valid_req_d ),
    .Q(\i_ibex/if_stage_i/prefetch_buffer_i/valid_req_q ),
    .Q_N(\i_ibex/if_stage_i/prefetch_buffer_i/valid_new_req_$_AND__A_B ),
    .CLK(clknet_leaf_149_clk_i_regs));
 sg13g2_buf_1 fanout437 (.A(\i_ibex/cs_registers_i/_0116_ ),
    .X(net437),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0494_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0069_ ),
    .B(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .A(\i_ibex/load_store_unit_i/ls_fsm_cs [2]));
 sg13g2_buf_2 fanout436 (.A(\i_ibex/cs_registers_i/_0116_ ),
    .X(net436),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout435 (.A(\i_ibex/ex_block_i/alu_adder_result_ext [2]),
    .X(net435),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0497_  (.A(net1461),
    .B(\i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ),
    .Y(\i_ibex/load_store_unit_i/_0072_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0498_  (.Y(\i_ibex/load_store_unit_i/_0073_ ),
    .B(\i_ibex/load_store_unit_i/_0072_ ),
    .A_N(net1462),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout434 (.X(net434),
    .A(net435),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0500_  (.Y(\i_ibex/load_store_unit_i/_0075_ ),
    .B(\i_ibex/load_store_unit_i/handle_misaligned_q ),
    .A_N(\i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg_E_$_AND__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0501_  (.Y(\i_ibex/lsu_addr_incr_req ),
    .B1(\i_ibex/load_store_unit_i/_0075_ ),
    .B2(net1462),
    .A2(\i_ibex/load_store_unit_i/_0073_ ),
    .A1(\i_ibex/load_store_unit_i/_0069_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout433 (.X(net433),
    .A(net434),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout432 (.A(net435),
    .X(net432),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/load_store_unit_i/_0504_  (.A(net688),
    .B_N(net471),
    .Y(\i_ibex/load_store_unit_i/_0078_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(net432),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/load_store_unit_i/_0506_  (.Y(\i_ibex/load_store_unit_i/_0080_ ),
    .A(\i_ibex/load_store_unit_i/pmp_err_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net432),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/load_store_unit_i/_0508_  (.A(net1757),
    .B_N(net1769),
    .Y(\i_ibex/load_store_unit_i/_0082_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/load_store_unit_i/_0509_  (.A(\i_ibex/load_store_unit_i/ls_fsm_cs [2]),
    .B(net1463),
    .C(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Y(\i_ibex/load_store_unit_i/_0083_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 \i_ibex/load_store_unit_i/_0510_  (.B(\i_ibex/load_store_unit_i/_0080_ ),
    .C(\i_ibex/load_store_unit_i/_0082_ ),
    .A(net1754),
    .Y(\i_ibex/load_store_unit_i/_0084_ ),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_ibex/load_store_unit_i/_0083_ ));
 sg13g2_nor3_2 \i_ibex/load_store_unit_i/_0511_  (.A(net1462),
    .B(net1460),
    .C(\i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ),
    .Y(\i_ibex/load_store_unit_i/_0085_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0512_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0086_ ),
    .A(\i_ibex/load_store_unit_i/lsu_err_q_$_NOT__A_Y ),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0513_  (.B1(net1460),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0087_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .A2(\i_ibex/load_store_unit_i/_0086_ ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0514_  (.A(net1754),
    .B(\i_ibex/load_store_unit_i/pmp_err_q ),
    .Y(\i_ibex/load_store_unit_i/_0088_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0515_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0089_ ),
    .B(\i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg_E_$_AND__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .A(net1459));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0516_  (.A(\i_ibex/load_store_unit_i/_0088_ ),
    .B(\i_ibex/load_store_unit_i/_0089_ ),
    .Y(\i_ibex/load_store_unit_i/_0090_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0517_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0091_ ),
    .A(net1459),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0518_  (.A(net1462),
    .B(net1460),
    .Y(\i_ibex/load_store_unit_i/_0092_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/load_store_unit_i/_0519_  (.A(net1754),
    .B(\i_ibex/lsu_req ),
    .X(\i_ibex/load_store_unit_i/_0093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/load_store_unit_i/_0520_  (.X(\i_ibex/load_store_unit_i/_0094_ ),
    .A(\i_ibex/load_store_unit_i/_0091_ ),
    .B(\i_ibex/load_store_unit_i/_0092_ ),
    .C(\i_ibex/load_store_unit_i/_0093_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0521_  (.VSS(VSS),
    .VDD(VDD),
    .B2(\i_ibex/load_store_unit_i/_0090_ ),
    .C1(\i_ibex/load_store_unit_i/_0094_ ),
    .B1(\i_ibex/load_store_unit_i/_0087_ ),
    .A1(\i_ibex/load_store_unit_i/_0082_ ),
    .Y(\i_ibex/load_store_unit_i/_0095_ ),
    .A2(\i_ibex/load_store_unit_i/_0085_ ));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0522_  (.VSS(VSS),
    .VDD(VDD),
    .B2(net1462),
    .C1(net1459),
    .B1(\i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg_E_$_AND__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .A1(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Y(\i_ibex/load_store_unit_i/_0096_ ),
    .A2(net1460));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0523_  (.A(\i_ibex/load_store_unit_i/_0085_ ),
    .B(\i_ibex/load_store_unit_i/_0096_ ),
    .Y(\i_ibex/load_store_unit_i/_0097_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/load_store_unit_i/_0524_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/load_store_unit_i/_0097_ ),
    .Y(\i_ibex/load_store_unit_i/_0098_ ),
    .A2(\i_ibex/load_store_unit_i/_0095_ ),
    .A1(\i_ibex/load_store_unit_i/_0084_ ));
 sg13g2_buf_4 fanout429 (.X(net429),
    .A(net432),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0526_  (.A0(\i_ibex/lsu_addr_last [0]),
    .A1(\i_ibex/load_store_unit_i/_0078_ ),
    .S(\i_ibex/load_store_unit_i/_0098_ ),
    .X(\i_ibex/load_store_unit_i/_0000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0527_  (.A0(\i_ibex/lsu_addr_last [10]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [11]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0001_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0528_  (.A0(\i_ibex/lsu_addr_last [11]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [12]),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0002_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0529_  (.A0(\i_ibex/lsu_addr_last [12]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [13]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0003_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0530_  (.A0(\i_ibex/lsu_addr_last [13]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [14]),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0004_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0531_  (.A0(\i_ibex/lsu_addr_last [14]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [15]),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0005_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0532_  (.A0(\i_ibex/lsu_addr_last [15]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [16]),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0533_  (.A0(\i_ibex/lsu_addr_last [16]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [17]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0007_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0534_  (.A0(\i_ibex/lsu_addr_last [17]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [18]),
    .S(net1136),
    .X(\i_ibex/load_store_unit_i/_0008_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0535_  (.A0(\i_ibex/lsu_addr_last [18]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [19]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0009_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(net432),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0537_  (.A0(\i_ibex/lsu_addr_last [19]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [20]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout427 (.A(\i_ibex/cs_registers_i/csr_wdata_int [20]),
    .X(net427),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/load_store_unit_i/_0540_  (.A(net688),
    .B_N(net433),
    .Y(\i_ibex/load_store_unit_i/_0103_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0541_  (.A0(\i_ibex/lsu_addr_last [1]),
    .A1(\i_ibex/load_store_unit_i/_0103_ ),
    .S(\i_ibex/load_store_unit_i/_0098_ ),
    .X(\i_ibex/load_store_unit_i/_0011_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0542_  (.A0(\i_ibex/lsu_addr_last [20]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [21]),
    .S(net1136),
    .X(\i_ibex/load_store_unit_i/_0012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0543_  (.A0(\i_ibex/lsu_addr_last [21]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [22]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0544_  (.A0(\i_ibex/lsu_addr_last [22]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [23]),
    .S(net1136),
    .X(\i_ibex/load_store_unit_i/_0014_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0545_  (.A0(\i_ibex/lsu_addr_last [23]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [24]),
    .S(net1136),
    .X(\i_ibex/load_store_unit_i/_0015_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0546_  (.A0(\i_ibex/lsu_addr_last [24]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [25]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0547_  (.A0(\i_ibex/lsu_addr_last [25]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [26]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0017_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0548_  (.A0(\i_ibex/lsu_addr_last [26]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [27]),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0549_  (.A0(\i_ibex/lsu_addr_last [27]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [28]),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0019_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout425 (.A(\i_ibex/cs_registers_i/csr_wdata_int [27]),
    .X(net425),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0551_  (.A0(\i_ibex/lsu_addr_last [28]),
    .A1(net1519),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0552_  (.A0(\i_ibex/lsu_addr_last [29]),
    .A1(net1518),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0553_  (.A0(\i_ibex/lsu_addr_last [2]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [3]),
    .S(net1137),
    .X(\i_ibex/load_store_unit_i/_0022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0554_  (.A0(\i_ibex/lsu_addr_last [30]),
    .A1(net1520),
    .S(net1135),
    .X(\i_ibex/load_store_unit_i/_0023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0555_  (.A0(\i_ibex/lsu_addr_last [31]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [32]),
    .S(net1136),
    .X(\i_ibex/load_store_unit_i/_0024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0556_  (.A0(\i_ibex/lsu_addr_last [3]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [4]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0025_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0557_  (.A0(\i_ibex/lsu_addr_last [4]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [5]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0558_  (.A0(\i_ibex/lsu_addr_last [5]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [6]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0027_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0559_  (.A0(\i_ibex/lsu_addr_last [6]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [7]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0560_  (.A0(\i_ibex/lsu_addr_last [7]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [8]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0561_  (.A0(\i_ibex/lsu_addr_last [8]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [9]),
    .S(net1133),
    .X(\i_ibex/load_store_unit_i/_0030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0562_  (.A0(\i_ibex/lsu_addr_last [9]),
    .A1(\i_ibex/ex_block_i/alu_adder_result_ext [10]),
    .S(net1134),
    .X(\i_ibex/load_store_unit_i/_0031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 \i_ibex/load_store_unit_i/_0563_  (.A(net1459),
    .B(net1463),
    .C(net1461),
    .Y(\i_ibex/load_store_unit_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/load_store_unit_i/_0564_  (.Y(\i_ibex/lsu_busy ),
    .A(\i_ibex/load_store_unit_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0566_  (.A(net1464),
    .B(\i_ibex/lsu_type [1]),
    .Y(\i_ibex/load_store_unit_i/_0107_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0567_  (.Y(\i_ibex/load_store_unit_i/_0108_ ),
    .B1(\i_ibex/load_store_unit_i/_0107_ ),
    .B2(\i_ibex/lsu_type [0]),
    .A2(\i_ibex/lsu_type [1]),
    .A1(net471),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0568_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0109_ ),
    .A(\i_ibex/load_store_unit_i/_0108_ ),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0569_  (.A(\i_ibex/lsu_type [0]),
    .B(\i_ibex/lsu_type [1]),
    .Y(\i_ibex/load_store_unit_i/_0110_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0570_  (.Y(\i_ibex/load_store_unit_i/_0111_ ),
    .B1(\i_ibex/load_store_unit_i/_0110_ ),
    .B2(\i_ibex/load_store_unit_i/data_be_o_$_MUX__Y_A [3]),
    .A2(\i_ibex/load_store_unit_i/_0109_ ),
    .A1(net433),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_16 \i_ibex/load_store_unit_i/_0571_  (.A(\i_ibex/load_store_unit_i/_0111_ ),
    .Y(data_be_o[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0572_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0112_ ),
    .A(\i_ibex/lsu_type [0]),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0573_  (.B(net1464),
    .C(\i_ibex/load_store_unit_i/_0112_ ),
    .A(net433),
    .Y(\i_ibex/load_store_unit_i/_0113_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0574_  (.B1(\i_ibex/load_store_unit_i/_0113_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0114_ ),
    .VSS(VSS),
    .A1(net433),
    .A2(net1464));
 sg13g2_nor3_1 \i_ibex/load_store_unit_i/_0575_  (.A(net471),
    .B(net1464),
    .C(\i_ibex/lsu_type [0]),
    .Y(\i_ibex/load_store_unit_i/_0115_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0576_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net471),
    .A2(\i_ibex/load_store_unit_i/_0114_ ),
    .Y(\i_ibex/load_store_unit_i/_0116_ ),
    .B1(\i_ibex/load_store_unit_i/_0115_ ));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0577_  (.Y(\i_ibex/load_store_unit_i/_0117_ ),
    .B(net1464),
    .A_N(\i_ibex/lsu_type [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/load_store_unit_i/_0578_  (.B(net434),
    .C(\i_ibex/load_store_unit_i/_0117_ ),
    .Y(\i_ibex/load_store_unit_i/_0118_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(net471));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0579_  (.B1(\i_ibex/load_store_unit_i/_0118_ ),
    .VDD(VDD),
    .Y(data_be_o[2]),
    .VSS(VSS),
    .A1(\i_ibex/lsu_type [1]),
    .A2(\i_ibex/load_store_unit_i/_0116_ ));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0580_  (.VSS(VSS),
    .VDD(VDD),
    .A1(net471),
    .A2(\i_ibex/lsu_type [1]),
    .Y(\i_ibex/load_store_unit_i/_0119_ ),
    .B1(\i_ibex/load_store_unit_i/_0107_ ));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0581_  (.B(net1464),
    .C(\i_ibex/load_store_unit_i/_0110_ ),
    .A(net434),
    .Y(\i_ibex/load_store_unit_i/_0120_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0582_  (.B1(\i_ibex/load_store_unit_i/_0120_ ),
    .VDD(VDD),
    .Y(data_be_o[1]),
    .VSS(VSS),
    .A1(net433),
    .A2(\i_ibex/load_store_unit_i/_0119_ ));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0583_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0121_ ),
    .B(net433),
    .A(net471));
 sg13g2_nor3_1 \i_ibex/load_store_unit_i/_0584_  (.A(\i_ibex/lsu_type [0]),
    .B(\i_ibex/load_store_unit_i/_0117_ ),
    .C(\i_ibex/load_store_unit_i/_0121_ ),
    .Y(\i_ibex/load_store_unit_i/_0122_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/load_store_unit_i/_0585_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/load_store_unit_i/_0122_ ),
    .Y(data_be_o[0]),
    .A2(\i_ibex/load_store_unit_i/_0121_ ),
    .A1(\i_ibex/load_store_unit_i/_0117_ ));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0586_  (.Y(\i_ibex/load_store_unit_i/_0123_ ),
    .A(\i_ibex/lsu_req ),
    .B(\i_ibex/load_store_unit_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/load_store_unit_i/_0587_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/load_store_unit_i/_0089_ ),
    .Y(\i_ibex/load_store_unit_i/_0124_ ),
    .A2(net1460),
    .A1(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0588_  (.A(\i_ibex/load_store_unit_i/_0083_ ),
    .B(\i_ibex/load_store_unit_i/_0124_ ),
    .Y(\i_ibex/load_store_unit_i/_0125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 \i_ibex/load_store_unit_i/_0589_  (.Y(data_req_o),
    .A(\i_ibex/load_store_unit_i/_0123_ ),
    .B(\i_ibex/load_store_unit_i/_0125_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0590_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0126_ ),
    .B(\i_ibex/load_store_unit_i/pmp_err_q ),
    .A(net1754));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0591_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0126_ ),
    .A2(\i_ibex/load_store_unit_i/_0124_ ),
    .Y(\i_ibex/load_store_unit_i/_0127_ ),
    .B1(\i_ibex/load_store_unit_i/_0094_ ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0592_  (.A(\i_ibex/load_store_unit_i/_0105_ ),
    .B(\i_ibex/load_store_unit_i/_0124_ ),
    .Y(\i_ibex/load_store_unit_i/_0128_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/load_store_unit_i/_0593_  (.A(\i_ibex/load_store_unit_i/_0127_ ),
    .B(\i_ibex/load_store_unit_i/_0128_ ),
    .Y(\i_ibex/load_store_unit_i/_0129_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0594_  (.A0(\i_ibex/load_store_unit_i/data_sign_ext_q ),
    .A1(\i_ibex/lsu_sign_ext ),
    .S(\i_ibex/load_store_unit_i/_0129_ ),
    .X(\i_ibex/load_store_unit_i/_0032_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0595_  (.A0(\i_ibex/load_store_unit_i/data_type_q [0]),
    .A1(\i_ibex/lsu_type [0]),
    .S(\i_ibex/load_store_unit_i/_0129_ ),
    .X(\i_ibex/load_store_unit_i/_0033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0596_  (.A0(\i_ibex/load_store_unit_i/data_type_q [1]),
    .A1(\i_ibex/lsu_type [1]),
    .S(\i_ibex/load_store_unit_i/_0129_ ),
    .X(\i_ibex/load_store_unit_i/_0034_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0597_  (.A0(\i_ibex/rf_rdata_b [31]),
    .A1(\i_ibex/rf_rdata_b [15]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0130_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0598_  (.A0(\i_ibex/rf_rdata_b [23]),
    .A1(\i_ibex/rf_rdata_b [7]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0131_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0600_  (.A0(\i_ibex/load_store_unit_i/_0130_ ),
    .A1(\i_ibex/load_store_unit_i/_0131_ ),
    .S(net468),
    .X(data_wdata_o[31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0602_  (.A0(\i_ibex/rf_rdata_b [30]),
    .A1(\i_ibex/rf_rdata_b [14]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0134_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0603_  (.A0(\i_ibex/rf_rdata_b [22]),
    .A1(\i_ibex/rf_rdata_b [6]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0135_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0604_  (.A0(\i_ibex/load_store_unit_i/_0134_ ),
    .A1(\i_ibex/load_store_unit_i/_0135_ ),
    .S(net468),
    .X(data_wdata_o[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0605_  (.A0(\i_ibex/rf_rdata_b [21]),
    .A1(\i_ibex/rf_rdata_b [5]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0136_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0606_  (.A0(\i_ibex/rf_rdata_b [13]),
    .A1(\i_ibex/rf_rdata_b [29]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0137_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0607_  (.A0(\i_ibex/load_store_unit_i/_0136_ ),
    .A1(\i_ibex/load_store_unit_i/_0137_ ),
    .S(net468),
    .X(data_wdata_o[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0608_  (.A0(\i_ibex/rf_rdata_b [20]),
    .A1(\i_ibex/rf_rdata_b [4]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0138_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0609_  (.A0(\i_ibex/rf_rdata_b [12]),
    .A1(\i_ibex/rf_rdata_b [28]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0139_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0610_  (.A0(\i_ibex/load_store_unit_i/_0138_ ),
    .A1(\i_ibex/load_store_unit_i/_0139_ ),
    .S(net468),
    .X(data_wdata_o[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0611_  (.A0(\i_ibex/rf_rdata_b [19]),
    .A1(\i_ibex/rf_rdata_b [3]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0140_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0612_  (.A0(\i_ibex/rf_rdata_b [11]),
    .A1(\i_ibex/rf_rdata_b [27]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0141_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0613_  (.A0(\i_ibex/load_store_unit_i/_0140_ ),
    .A1(\i_ibex/load_store_unit_i/_0141_ ),
    .S(net467),
    .X(data_wdata_o[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0614_  (.A0(\i_ibex/rf_rdata_b [18]),
    .A1(\i_ibex/rf_rdata_b [2]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0142_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0615_  (.A0(\i_ibex/rf_rdata_b [10]),
    .A1(\i_ibex/rf_rdata_b [26]),
    .S(net428),
    .X(\i_ibex/load_store_unit_i/_0143_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0616_  (.A0(\i_ibex/load_store_unit_i/_0142_ ),
    .A1(\i_ibex/load_store_unit_i/_0143_ ),
    .S(net467),
    .X(data_wdata_o[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout421 (.A(\i_ibex/cs_registers_i/csr_wdata_int [29]),
    .X(net421),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0618_  (.A0(\i_ibex/rf_rdata_b [17]),
    .A1(\i_ibex/rf_rdata_b [1]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0145_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0619_  (.A0(\i_ibex/rf_rdata_b [9]),
    .A1(\i_ibex/rf_rdata_b [25]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0146_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0620_  (.A0(\i_ibex/load_store_unit_i/_0145_ ),
    .A1(\i_ibex/load_store_unit_i/_0146_ ),
    .S(net467),
    .X(data_wdata_o[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0621_  (.A0(\i_ibex/rf_rdata_b [16]),
    .A1(net1513),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0147_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0622_  (.A0(\i_ibex/rf_rdata_b [8]),
    .A1(\i_ibex/rf_rdata_b [24]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0148_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0623_  (.A0(\i_ibex/load_store_unit_i/_0147_ ),
    .A1(\i_ibex/load_store_unit_i/_0148_ ),
    .S(net467),
    .X(data_wdata_o[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0624_  (.A0(\i_ibex/rf_rdata_b [15]),
    .A1(\i_ibex/rf_rdata_b [31]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0149_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0625_  (.A0(\i_ibex/rf_rdata_b [7]),
    .A1(\i_ibex/rf_rdata_b [23]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0150_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0626_  (.A0(\i_ibex/load_store_unit_i/_0149_ ),
    .A1(\i_ibex/load_store_unit_i/_0150_ ),
    .S(net467),
    .X(data_wdata_o[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0627_  (.A0(\i_ibex/rf_rdata_b [14]),
    .A1(\i_ibex/rf_rdata_b [30]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0151_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0628_  (.A0(\i_ibex/rf_rdata_b [6]),
    .A1(\i_ibex/rf_rdata_b [22]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0152_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0630_  (.A0(\i_ibex/load_store_unit_i/_0151_ ),
    .A1(\i_ibex/load_store_unit_i/_0152_ ),
    .S(net469),
    .X(data_wdata_o[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0631_  (.A0(\i_ibex/rf_rdata_b [5]),
    .A1(\i_ibex/rf_rdata_b [21]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0154_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0632_  (.A0(\i_ibex/load_store_unit_i/_0137_ ),
    .A1(\i_ibex/load_store_unit_i/_0154_ ),
    .S(net469),
    .X(data_wdata_o[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0633_  (.A0(\i_ibex/rf_rdata_b [4]),
    .A1(\i_ibex/rf_rdata_b [20]),
    .S(net429),
    .X(\i_ibex/load_store_unit_i/_0155_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0634_  (.A0(\i_ibex/load_store_unit_i/_0139_ ),
    .A1(\i_ibex/load_store_unit_i/_0155_ ),
    .S(net469),
    .X(data_wdata_o[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0636_  (.A0(\i_ibex/rf_rdata_b [29]),
    .A1(\i_ibex/rf_rdata_b [13]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0157_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0637_  (.A0(\i_ibex/load_store_unit_i/_0157_ ),
    .A1(\i_ibex/load_store_unit_i/_0136_ ),
    .S(net469),
    .X(data_wdata_o[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0638_  (.A0(\i_ibex/rf_rdata_b [3]),
    .A1(\i_ibex/rf_rdata_b [19]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0158_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0639_  (.A0(\i_ibex/load_store_unit_i/_0141_ ),
    .A1(\i_ibex/load_store_unit_i/_0158_ ),
    .S(net469),
    .X(data_wdata_o[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0640_  (.A0(\i_ibex/rf_rdata_b [2]),
    .A1(\i_ibex/rf_rdata_b [18]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0159_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0641_  (.A0(\i_ibex/load_store_unit_i/_0143_ ),
    .A1(\i_ibex/load_store_unit_i/_0159_ ),
    .S(net469),
    .X(data_wdata_o[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0642_  (.A0(\i_ibex/rf_rdata_b [1]),
    .A1(\i_ibex/rf_rdata_b [17]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0160_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0643_  (.A0(\i_ibex/load_store_unit_i/_0146_ ),
    .A1(\i_ibex/load_store_unit_i/_0160_ ),
    .S(net468),
    .X(data_wdata_o[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0644_  (.A0(net1513),
    .A1(\i_ibex/rf_rdata_b [16]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0161_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0645_  (.A0(\i_ibex/load_store_unit_i/_0148_ ),
    .A1(\i_ibex/load_store_unit_i/_0161_ ),
    .S(net468),
    .X(data_wdata_o[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0646_  (.A0(\i_ibex/load_store_unit_i/_0150_ ),
    .A1(\i_ibex/load_store_unit_i/_0130_ ),
    .S(net468),
    .X(data_wdata_o[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0647_  (.A0(\i_ibex/load_store_unit_i/_0152_ ),
    .A1(\i_ibex/load_store_unit_i/_0134_ ),
    .S(net468),
    .X(data_wdata_o[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0649_  (.A0(\i_ibex/load_store_unit_i/_0154_ ),
    .A1(\i_ibex/load_store_unit_i/_0157_ ),
    .S(net470),
    .X(data_wdata_o[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0650_  (.A0(\i_ibex/rf_rdata_b [28]),
    .A1(\i_ibex/rf_rdata_b [12]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0163_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0651_  (.A0(\i_ibex/load_store_unit_i/_0155_ ),
    .A1(\i_ibex/load_store_unit_i/_0163_ ),
    .S(net470),
    .X(data_wdata_o[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0652_  (.A0(\i_ibex/rf_rdata_b [27]),
    .A1(\i_ibex/rf_rdata_b [11]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0164_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0653_  (.A0(\i_ibex/load_store_unit_i/_0158_ ),
    .A1(\i_ibex/load_store_unit_i/_0164_ ),
    .S(net470),
    .X(data_wdata_o[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0654_  (.A0(\i_ibex/rf_rdata_b [26]),
    .A1(\i_ibex/rf_rdata_b [10]),
    .S(net431),
    .X(\i_ibex/load_store_unit_i/_0165_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0655_  (.A0(\i_ibex/load_store_unit_i/_0159_ ),
    .A1(\i_ibex/load_store_unit_i/_0165_ ),
    .S(net470),
    .X(data_wdata_o[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0656_  (.A0(\i_ibex/load_store_unit_i/_0163_ ),
    .A1(\i_ibex/load_store_unit_i/_0138_ ),
    .S(net470),
    .X(data_wdata_o[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0657_  (.A0(\i_ibex/rf_rdata_b [25]),
    .A1(\i_ibex/rf_rdata_b [9]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0166_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0658_  (.A0(\i_ibex/load_store_unit_i/_0160_ ),
    .A1(\i_ibex/load_store_unit_i/_0166_ ),
    .S(net470),
    .X(data_wdata_o[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0659_  (.A0(\i_ibex/rf_rdata_b [24]),
    .A1(\i_ibex/rf_rdata_b [8]),
    .S(net430),
    .X(\i_ibex/load_store_unit_i/_0167_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0660_  (.A0(\i_ibex/load_store_unit_i/_0161_ ),
    .A1(\i_ibex/load_store_unit_i/_0167_ ),
    .S(net470),
    .X(data_wdata_o[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0661_  (.A0(\i_ibex/load_store_unit_i/_0164_ ),
    .A1(\i_ibex/load_store_unit_i/_0140_ ),
    .S(net470),
    .X(data_wdata_o[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0662_  (.A0(\i_ibex/load_store_unit_i/_0165_ ),
    .A1(\i_ibex/load_store_unit_i/_0142_ ),
    .S(net469),
    .X(data_wdata_o[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0663_  (.A0(\i_ibex/load_store_unit_i/_0166_ ),
    .A1(\i_ibex/load_store_unit_i/_0145_ ),
    .S(net469),
    .X(data_wdata_o[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0664_  (.A0(\i_ibex/load_store_unit_i/_0167_ ),
    .A1(\i_ibex/load_store_unit_i/_0147_ ),
    .S(net467),
    .X(data_wdata_o[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0665_  (.A0(\i_ibex/load_store_unit_i/_0131_ ),
    .A1(\i_ibex/load_store_unit_i/_0149_ ),
    .S(net467),
    .X(data_wdata_o[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_2 \i_ibex/load_store_unit_i/_0666_  (.A0(\i_ibex/load_store_unit_i/_0135_ ),
    .A1(\i_ibex/load_store_unit_i/_0151_ ),
    .S(net467),
    .X(data_wdata_o[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0667_  (.A0(\i_ibex/load_store_unit_i/data_we_q ),
    .A1(\i_ibex/lsu_we ),
    .S(\i_ibex/load_store_unit_i/_0129_ ),
    .X(\i_ibex/load_store_unit_i/_0035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/load_store_unit_i/_0668_  (.A(net1769),
    .B(\i_ibex/load_store_unit_i/pmp_err_q ),
    .Y(\i_ibex/load_store_unit_i/_0168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/load_store_unit_i/_0669_  (.A(net1754),
    .B(net1463),
    .C(\i_ibex/load_store_unit_i/_0069_ ),
    .D(\i_ibex/load_store_unit_i/_0168_ ),
    .Y(\i_ibex/load_store_unit_i/_0169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0670_  (.A(net1460),
    .B(\i_ibex/load_store_unit_i/_0089_ ),
    .Y(\i_ibex/load_store_unit_i/_0170_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0671_  (.B1(\i_ibex/load_store_unit_i/_0170_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0171_ ),
    .VSS(VSS),
    .A1(net1464),
    .A2(\i_ibex/load_store_unit_i/_0126_ ));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0672_  (.Y(\i_ibex/load_store_unit_i/_0172_ ),
    .B(\i_ibex/load_store_unit_i/_0171_ ),
    .A_N(\i_ibex/load_store_unit_i/_0169_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0673_  (.B1(net471),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0173_ ),
    .VSS(VSS),
    .A1(net433),
    .A2(\i_ibex/load_store_unit_i/_0112_ ));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0674_  (.Y(\i_ibex/load_store_unit_i/_0174_ ),
    .A(net433),
    .B(\i_ibex/load_store_unit_i/_0112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0675_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0173_ ),
    .A2(\i_ibex/load_store_unit_i/_0174_ ),
    .Y(\i_ibex/load_store_unit_i/_0175_ ),
    .B1(\i_ibex/lsu_type [1]));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0676_  (.A0(\i_ibex/load_store_unit_i/_0172_ ),
    .A1(\i_ibex/load_store_unit_i/_0175_ ),
    .S(\i_ibex/load_store_unit_i/_0125_ ),
    .X(\i_ibex/load_store_unit_i/_0176_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0677_  (.B1(\i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg_E_$_AND__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0177_ ),
    .VSS(VSS),
    .A1(net1463),
    .A2(net1769));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0678_  (.A(\i_ibex/load_store_unit_i/_0069_ ),
    .B(\i_ibex/load_store_unit_i/_0126_ ),
    .Y(\i_ibex/load_store_unit_i/_0178_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0679_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0177_ ),
    .A2(\i_ibex/load_store_unit_i/_0178_ ),
    .Y(\i_ibex/load_store_unit_i/_0179_ ),
    .B1(\i_ibex/load_store_unit_i/_0105_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0680_  (.B1(\i_ibex/load_store_unit_i/_0096_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0180_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0093_ ),
    .A2(\i_ibex/load_store_unit_i/_0179_ ));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0681_  (.A0(\i_ibex/load_store_unit_i/_0176_ ),
    .A1(net1464),
    .S(\i_ibex/load_store_unit_i/_0180_ ),
    .X(\i_ibex/load_store_unit_i/_0036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/load_store_unit_i/_0682_  (.A(\i_ibex/lsu_busy ),
    .B(\i_ibex/load_store_unit_i/_0168_ ),
    .Y(\i_ibex/lsu_resp_valid ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0683_  (.B1(net1769),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0181_ ),
    .VSS(VSS),
    .A1(net1757),
    .A2(\i_ibex/load_store_unit_i/lsu_err_q ));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0684_  (.Y(\i_ibex/load_store_unit_i/_0182_ ),
    .A(\i_ibex/load_store_unit_i/lsu_rdata_valid_o_$_AND__Y_B ),
    .B(\i_ibex/load_store_unit_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/load_store_unit_i/_0685_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/load_store_unit_i/_0182_ ),
    .Y(\i_ibex/lsu_load_err ),
    .A2(\i_ibex/load_store_unit_i/_0181_ ),
    .A1(\i_ibex/load_store_unit_i/_0080_ ));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0686_  (.Y(\i_ibex/load_store_unit_i/_0183_ ),
    .B(\i_ibex/load_store_unit_i/_0083_ ),
    .A_N(\i_ibex/load_store_unit_i/_0168_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0687_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/lsu_busy ),
    .A2(\i_ibex/load_store_unit_i/_0183_ ),
    .Y(\i_ibex/load_store_unit_i/_0184_ ),
    .B1(net1754));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0688_  (.A(net1459),
    .B(\i_ibex/lsu_req ),
    .Y(\i_ibex/load_store_unit_i/_0185_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0689_  (.A(\i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ),
    .B(net1769),
    .Y(\i_ibex/load_store_unit_i/_0186_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0690_  (.B1(\i_ibex/load_store_unit_i/_0092_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0187_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0185_ ),
    .A2(\i_ibex/load_store_unit_i/_0186_ ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0691_  (.A(net1459),
    .B(net1462),
    .Y(\i_ibex/load_store_unit_i/_0188_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0692_  (.Y(\i_ibex/load_store_unit_i/_0189_ ),
    .B(\i_ibex/load_store_unit_i/_0188_ ),
    .A_N(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0693_  (.A(net1769),
    .B(\i_ibex/load_store_unit_i/_0189_ ),
    .Y(\i_ibex/load_store_unit_i/_0190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0694_  (.B1(\i_ibex/load_store_unit_i/_0088_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0191_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0124_ ),
    .A2(\i_ibex/load_store_unit_i/_0190_ ));
 sg13g2_nand2_2 \i_ibex/load_store_unit_i/_0695_  (.Y(\i_ibex/load_store_unit_i/_0192_ ),
    .A(\i_ibex/load_store_unit_i/_0187_ ),
    .B(\i_ibex/load_store_unit_i/_0191_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0696_  (.A0(net1755),
    .A1(net1463),
    .S(\i_ibex/load_store_unit_i/_0192_ ),
    .X(\i_ibex/load_store_unit_i/_0037_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 \i_ibex/load_store_unit_i/_0697_  (.B(\i_ibex/load_store_unit_i/_0175_ ),
    .A(net1754),
    .X(\i_ibex/load_store_unit_i/_0193_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0698_  (.A(\i_ibex/load_store_unit_i/_0169_ ),
    .B(\i_ibex/load_store_unit_i/_0170_ ),
    .Y(\i_ibex/load_store_unit_i/_0194_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0699_  (.B1(\i_ibex/load_store_unit_i/_0194_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0195_ ),
    .VSS(VSS),
    .A1(\i_ibex/lsu_busy ),
    .A2(\i_ibex/load_store_unit_i/_0193_ ));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0700_  (.A0(\i_ibex/load_store_unit_i/_0195_ ),
    .A1(net1460),
    .S(\i_ibex/load_store_unit_i/_0192_ ),
    .X(\i_ibex/load_store_unit_i/_0038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 \i_ibex/load_store_unit_i/_0701_  (.A(\i_ibex/load_store_unit_i/_0083_ ),
    .B(\i_ibex/load_store_unit_i/_0168_ ),
    .X(\i_ibex/load_store_unit_i/_0196_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0702_  (.A0(\i_ibex/load_store_unit_i/_0196_ ),
    .A1(net1459),
    .S(\i_ibex/load_store_unit_i/_0192_ ),
    .X(\i_ibex/load_store_unit_i/_0039_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0703_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0197_ ),
    .B(\i_ibex/load_store_unit_i/pmp_err_q ),
    .A(net1757));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0704_  (.Y(\i_ibex/load_store_unit_i/_0198_ ),
    .B1(\i_ibex/load_store_unit_i/_0083_ ),
    .B2(\i_ibex/load_store_unit_i/_0197_ ),
    .A2(\i_ibex/load_store_unit_i/_0085_ ),
    .A1(net1757),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0705_  (.A(\i_ibex/load_store_unit_i/_0091_ ),
    .B(\i_ibex/load_store_unit_i/_0072_ ),
    .Y(\i_ibex/load_store_unit_i/_0199_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/load_store_unit_i/_0706_  (.A(net1461),
    .B_N(\i_ibex/lsu_req ),
    .Y(\i_ibex/load_store_unit_i/_0200_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/load_store_unit_i/_0707_  (.A(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .B_N(net1461),
    .Y(\i_ibex/load_store_unit_i/_0201_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 \i_ibex/load_store_unit_i/_0708_  (.A(net1459),
    .B(\i_ibex/load_store_unit_i/_0200_ ),
    .C(\i_ibex/load_store_unit_i/_0201_ ),
    .Y(\i_ibex/load_store_unit_i/_0202_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0709_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0080_ ),
    .A2(\i_ibex/load_store_unit_i/_0083_ ),
    .Y(\i_ibex/load_store_unit_i/_0203_ ),
    .B1(\i_ibex/load_store_unit_i/_0085_ ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0710_  (.A(data_rvalid_i),
    .B(\i_ibex/load_store_unit_i/_0203_ ),
    .Y(\i_ibex/load_store_unit_i/_0204_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/load_store_unit_i/_0711_  (.A(net1462),
    .B(\i_ibex/load_store_unit_i/_0199_ ),
    .C(\i_ibex/load_store_unit_i/_0202_ ),
    .D(\i_ibex/load_store_unit_i/_0204_ ),
    .Y(\i_ibex/load_store_unit_i/_0205_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0712_  (.A(\i_ibex/load_store_unit_i/lsu_err_q ),
    .B(\i_ibex/load_store_unit_i/_0205_ ),
    .Y(\i_ibex/load_store_unit_i/_0206_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0713_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0198_ ),
    .A2(\i_ibex/load_store_unit_i/_0205_ ),
    .Y(\i_ibex/load_store_unit_i/_0040_ ),
    .B1(\i_ibex/load_store_unit_i/_0206_ ));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0714_  (.A2(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_1_Y ),
    .A1(\i_ibex/load_store_unit_i/data_type_q [1]),
    .B1(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_Y ),
    .X(\i_ibex/load_store_unit_i/_0207_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0715_  (.B1(\i_ibex/load_store_unit_i/_0207_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0208_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/data_type_q [0]),
    .A2(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_1_Y ));
 sg13g2_buf_2 fanout417 (.A(\i_ibex/cs_registers_i/csr_wdata_int [25]),
    .X(net417),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0718_  (.A(\i_ibex/load_store_unit_i/rdata_offset_q [0]),
    .B(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_1_Y ),
    .Y(\i_ibex/load_store_unit_i/_0211_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout415 (.A(\i_ibex/cs_registers_i/csr_wdata_int [23]),
    .X(net415),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout413 (.A(\i_ibex/cs_registers_i/csr_wdata_int [22]),
    .X(net413),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0722_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/rdata_offset_q [1]),
    .A2(net1458),
    .Y(\i_ibex/load_store_unit_i/_0215_ ),
    .B1(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0723_  (.A(net1428),
    .B(\i_ibex/load_store_unit_i/_0215_ ),
    .Y(\i_ibex/load_store_unit_i/_0216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(\i_ibex/cs_registers_i/csr_wdata_int [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout411 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_099_ ),
    .X(net411),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0726_  (.A(\i_ibex/load_store_unit_i/rdata_offset_q [1]),
    .B(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .Y(\i_ibex/load_store_unit_i/_0219_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout410 (.A(\i_ibex/cs_registers_i/minstret_counter_i_counter_inc_i ),
    .X(net410),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout409 (.A(\i_ibex/cs_registers_i/minstret_counter_i_counter_inc_i ),
    .X(net409),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0729_  (.A(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .B(net1458),
    .Y(\i_ibex/load_store_unit_i/_0222_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout408 (.A(\i_ibex/cs_registers_i/minstret_counter_i_counter_inc_i ),
    .X(net408),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout407 (.A(\i_ibex/cs_registers_i/mhpmcounterh_we [0]),
    .X(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0732_  (.Y(\i_ibex/load_store_unit_i/_0225_ ),
    .B1(net1412),
    .B2(data_rdata_i[23]),
    .A2(net1418),
    .A1(data_rdata_i[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0733_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0226_ ),
    .A(\i_ibex/load_store_unit_i/_0225_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0734_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[31]),
    .C1(\i_ibex/load_store_unit_i/_0226_ ),
    .B1(net1403),
    .A1(data_rdata_i[15]),
    .Y(\i_ibex/load_store_unit_i/_0227_ ),
    .A2(net1429));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0735_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0228_ ),
    .A(net1458),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0736_  (.Y(\i_ibex/load_store_unit_i/_0229_ ),
    .A(\i_ibex/load_store_unit_i/rdata_offset_q [0]),
    .B(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0737_  (.B1(\i_ibex/load_store_unit_i/_0229_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0230_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0228_ ),
    .A2(net1418));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0738_  (.Y(\i_ibex/load_store_unit_i/_0231_ ),
    .B(data_rdata_i[31]),
    .A_N(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0739_  (.Y(\i_ibex/load_store_unit_i/_0232_ ),
    .B(data_rdata_i[23]),
    .A_N(\i_ibex/load_store_unit_i/rdata_offset_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0740_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0231_ ),
    .A2(\i_ibex/load_store_unit_i/_0232_ ),
    .Y(\i_ibex/load_store_unit_i/_0233_ ),
    .B1(net1458));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0741_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[7]),
    .C1(\i_ibex/load_store_unit_i/_0233_ ),
    .B1(\i_ibex/load_store_unit_i/_0230_ ),
    .A1(data_rdata_i[15]),
    .Y(\i_ibex/load_store_unit_i/_0234_ ),
    .A2(net1419));
 sg13g2_a21oi_2 \i_ibex/load_store_unit_i/_0742_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_1_Y ),
    .Y(\i_ibex/load_store_unit_i/_0235_ ),
    .A2(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_Y ),
    .A1(\i_ibex/load_store_unit_i/data_type_q [0]));
 sg13g2_nand3b_1 \i_ibex/load_store_unit_i/_0743_  (.B(net1457),
    .C(\i_ibex/load_store_unit_i/data_sign_ext_q ),
    .Y(\i_ibex/load_store_unit_i/_0236_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/load_store_unit_i/_0234_ ));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0745_  (.Y(\i_ibex/load_store_unit_i/_0238_ ),
    .B(data_rdata_i[7]),
    .A_N(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0746_  (.Y(\i_ibex/load_store_unit_i/_0239_ ),
    .B(data_rdata_i[31]),
    .A_N(\i_ibex/load_store_unit_i/rdata_offset_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0747_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0238_ ),
    .A2(\i_ibex/load_store_unit_i/_0239_ ),
    .Y(\i_ibex/load_store_unit_i/_0240_ ),
    .B1(net1458));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0748_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[15]),
    .C1(\i_ibex/load_store_unit_i/_0240_ ),
    .B1(\i_ibex/load_store_unit_i/_0230_ ),
    .A1(data_rdata_i[23]),
    .Y(\i_ibex/load_store_unit_i/_0241_ ),
    .A2(net1419));
 sg13g2_nor2_2 \i_ibex/load_store_unit_i/_0749_  (.A(\i_ibex/load_store_unit_i/data_type_q [1]),
    .B(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_Y ),
    .Y(\i_ibex/load_store_unit_i/_0242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 \i_ibex/load_store_unit_i/_0750_  (.B(net1456),
    .C(\i_ibex/load_store_unit_i/data_sign_ext_q ),
    .Y(\i_ibex/load_store_unit_i/_0243_ ),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\i_ibex/load_store_unit_i/_0241_ ));
 sg13g2_and2_1 \i_ibex/load_store_unit_i/_0751_  (.A(net635),
    .B(\i_ibex/load_store_unit_i/_0243_ ),
    .X(\i_ibex/load_store_unit_i/_0244_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(\i_ibex/cs_registers_i/mhpmcounterh_we [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0753_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [31]),
    .VSS(VSS),
    .A1(net1434),
    .A2(\i_ibex/load_store_unit_i/_0227_ ));
 sg13g2_buf_2 fanout404 (.A(net407),
    .X(net404),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0757_  (.Y(\i_ibex/load_store_unit_i/_0249_ ),
    .B1(net1409),
    .B2(data_rdata_i[22]),
    .A2(net1423),
    .A1(data_rdata_i[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0758_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0250_ ),
    .A(\i_ibex/load_store_unit_i/_0249_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0759_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[30]),
    .C1(\i_ibex/load_store_unit_i/_0250_ ),
    .B1(net1400),
    .A1(data_rdata_i[6]),
    .Y(\i_ibex/load_store_unit_i/_0251_ ),
    .A2(net1414));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0760_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [30]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0251_ ));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0762_  (.Y(\i_ibex/load_store_unit_i/_0253_ ),
    .B1(net1410),
    .B2(data_rdata_i[13]),
    .A2(net1417),
    .A1(\i_ibex/load_store_unit_i/rdata_q [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0763_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0254_ ),
    .A(\i_ibex/load_store_unit_i/_0253_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0764_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[21]),
    .C1(\i_ibex/load_store_unit_i/_0254_ ),
    .B1(net1402),
    .A1(data_rdata_i[5]),
    .Y(\i_ibex/load_store_unit_i/_0255_ ),
    .A2(net1430));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0765_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [21]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0255_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0766_  (.Y(\i_ibex/load_store_unit_i/_0256_ ),
    .B1(net1411),
    .B2(data_rdata_i[12]),
    .A2(net1415),
    .A1(\i_ibex/load_store_unit_i/rdata_q [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0767_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0257_ ),
    .A(\i_ibex/load_store_unit_i/_0256_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0768_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[20]),
    .C1(\i_ibex/load_store_unit_i/_0257_ ),
    .B1(net1400),
    .A1(data_rdata_i[4]),
    .Y(\i_ibex/load_store_unit_i/_0258_ ),
    .A2(net1424));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0769_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [20]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0258_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0770_  (.Y(\i_ibex/load_store_unit_i/_0259_ ),
    .B1(net1410),
    .B2(data_rdata_i[11]),
    .A2(net1416),
    .A1(\i_ibex/load_store_unit_i/rdata_q [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0771_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0260_ ),
    .A(\i_ibex/load_store_unit_i/_0259_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0772_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[19]),
    .C1(\i_ibex/load_store_unit_i/_0260_ ),
    .B1(net1401),
    .A1(data_rdata_i[3]),
    .Y(\i_ibex/load_store_unit_i/_0261_ ),
    .A2(net1425));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0773_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [19]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0261_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0774_  (.Y(\i_ibex/load_store_unit_i/_0262_ ),
    .B1(net1413),
    .B2(data_rdata_i[10]),
    .A2(net1418),
    .A1(\i_ibex/load_store_unit_i/rdata_q [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0775_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0263_ ),
    .A(\i_ibex/load_store_unit_i/_0262_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0776_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[18]),
    .C1(\i_ibex/load_store_unit_i/_0263_ ),
    .B1(net1403),
    .A1(data_rdata_i[2]),
    .Y(\i_ibex/load_store_unit_i/_0264_ ),
    .A2(net1428));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0777_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [18]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0264_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0778_  (.Y(\i_ibex/load_store_unit_i/_0265_ ),
    .B1(net1409),
    .B2(data_rdata_i[9]),
    .A2(net1414),
    .A1(\i_ibex/load_store_unit_i/rdata_q [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0779_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0266_ ),
    .A(\i_ibex/load_store_unit_i/_0265_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0780_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[17]),
    .C1(\i_ibex/load_store_unit_i/_0266_ ),
    .B1(net1400),
    .A1(data_rdata_i[1]),
    .Y(\i_ibex/load_store_unit_i/_0267_ ),
    .A2(net1424));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0781_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [17]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0267_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0782_  (.Y(\i_ibex/load_store_unit_i/_0268_ ),
    .B1(net1413),
    .B2(data_rdata_i[8]),
    .A2(net1421),
    .A1(\i_ibex/load_store_unit_i/rdata_q [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0783_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0269_ ),
    .A(\i_ibex/load_store_unit_i/_0268_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0784_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[16]),
    .C1(\i_ibex/load_store_unit_i/_0269_ ),
    .B1(net1402),
    .A1(data_rdata_i[0]),
    .Y(\i_ibex/load_store_unit_i/_0270_ ),
    .A2(net1430));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0785_  (.B1(\i_ibex/load_store_unit_i/_0244_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [16]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0270_ ));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0787_  (.Y(\i_ibex/load_store_unit_i/_0272_ ),
    .B1(\i_ibex/load_store_unit_i/_0230_ ),
    .B2(data_rdata_i[15]),
    .A2(net1412),
    .A1(data_rdata_i[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0788_  (.Y(\i_ibex/load_store_unit_i/_0273_ ),
    .B1(net1429),
    .B2(data_rdata_i[31]),
    .A2(net1419),
    .A1(data_rdata_i[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 \i_ibex/load_store_unit_i/_0789_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0274_ ),
    .B(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_Y ),
    .A(\i_ibex/load_store_unit_i/data_type_q [1]));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0790_  (.A2(\i_ibex/load_store_unit_i/_0273_ ),
    .A1(\i_ibex/load_store_unit_i/_0272_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0275_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(net407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0793_  (.Y(\i_ibex/load_store_unit_i/_0278_ ),
    .B1(net1429),
    .B2(\i_ibex/load_store_unit_i/rdata_q [23]),
    .A2(net1419),
    .A1(\i_ibex/load_store_unit_i/rdata_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout397 (.A(\i_ibex/cs_registers_i/mcycle_counter_i/_091_ ),
    .X(net397),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0795_  (.A2(\i_ibex/load_store_unit_i/_0278_ ),
    .A1(\i_ibex/load_store_unit_i/_0272_ ),
    .B1(net1434),
    .X(\i_ibex/load_store_unit_i/_0280_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0796_  (.B(\i_ibex/load_store_unit_i/_0275_ ),
    .C(\i_ibex/load_store_unit_i/_0280_ ),
    .A(\i_ibex/load_store_unit_i/_0236_ ),
    .Y(\i_ibex/rf_wdata_lsu [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout396 (.A(net397),
    .X(net396),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0798_  (.Y(\i_ibex/load_store_unit_i/_0282_ ),
    .B1(net1400),
    .B2(data_rdata_i[14]),
    .A2(net1409),
    .A1(data_rdata_i[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0799_  (.Y(\i_ibex/load_store_unit_i/_0283_ ),
    .B1(net1423),
    .B2(data_rdata_i[30]),
    .A2(net1414),
    .A1(data_rdata_i[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0800_  (.A2(\i_ibex/load_store_unit_i/_0283_ ),
    .A1(\i_ibex/load_store_unit_i/_0282_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0284_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0801_  (.Y(\i_ibex/load_store_unit_i/_0285_ ),
    .B1(net1423),
    .B2(\i_ibex/load_store_unit_i/rdata_q [22]),
    .A2(net1414),
    .A1(\i_ibex/load_store_unit_i/rdata_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0802_  (.A2(\i_ibex/load_store_unit_i/_0285_ ),
    .A1(\i_ibex/load_store_unit_i/_0282_ ),
    .B1(net1432),
    .X(\i_ibex/load_store_unit_i/_0286_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0803_  (.B(\i_ibex/load_store_unit_i/_0284_ ),
    .C(\i_ibex/load_store_unit_i/_0286_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0804_  (.Y(\i_ibex/load_store_unit_i/_0287_ ),
    .B1(net1401),
    .B2(data_rdata_i[13]),
    .A2(net1411),
    .A1(data_rdata_i[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0805_  (.Y(\i_ibex/load_store_unit_i/_0288_ ),
    .B1(net1426),
    .B2(data_rdata_i[29]),
    .A2(net1417),
    .A1(data_rdata_i[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0806_  (.A2(\i_ibex/load_store_unit_i/_0288_ ),
    .A1(\i_ibex/load_store_unit_i/_0287_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0289_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0807_  (.Y(\i_ibex/load_store_unit_i/_0290_ ),
    .B1(net1426),
    .B2(\i_ibex/load_store_unit_i/rdata_q [21]),
    .A2(net1417),
    .A1(\i_ibex/load_store_unit_i/rdata_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0808_  (.A2(\i_ibex/load_store_unit_i/_0290_ ),
    .A1(\i_ibex/load_store_unit_i/_0287_ ),
    .B1(net1436),
    .X(\i_ibex/load_store_unit_i/_0291_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0809_  (.B(\i_ibex/load_store_unit_i/_0289_ ),
    .C(\i_ibex/load_store_unit_i/_0291_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0810_  (.Y(\i_ibex/load_store_unit_i/_0292_ ),
    .B1(net1403),
    .B2(data_rdata_i[12]),
    .A2(net1412),
    .A1(data_rdata_i[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0811_  (.Y(\i_ibex/load_store_unit_i/_0293_ ),
    .B1(net1428),
    .B2(data_rdata_i[28]),
    .A2(net1418),
    .A1(data_rdata_i[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0812_  (.A2(\i_ibex/load_store_unit_i/_0293_ ),
    .A1(\i_ibex/load_store_unit_i/_0292_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0294_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0813_  (.Y(\i_ibex/load_store_unit_i/_0295_ ),
    .B1(net1428),
    .B2(\i_ibex/load_store_unit_i/rdata_q [20]),
    .A2(net1418),
    .A1(\i_ibex/load_store_unit_i/rdata_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0814_  (.A2(\i_ibex/load_store_unit_i/_0295_ ),
    .A1(\i_ibex/load_store_unit_i/_0292_ ),
    .B1(net1433),
    .X(\i_ibex/load_store_unit_i/_0296_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0815_  (.B(\i_ibex/load_store_unit_i/_0294_ ),
    .C(\i_ibex/load_store_unit_i/_0296_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0816_  (.Y(\i_ibex/load_store_unit_i/_0297_ ),
    .B1(net1410),
    .B2(data_rdata_i[21]),
    .A2(net1426),
    .A1(data_rdata_i[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0817_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0298_ ),
    .A(\i_ibex/load_store_unit_i/_0297_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0818_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[29]),
    .C1(\i_ibex/load_store_unit_i/_0298_ ),
    .B1(net1402),
    .A1(data_rdata_i[5]),
    .Y(\i_ibex/load_store_unit_i/_0299_ ),
    .A2(net1420));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0819_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [29]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0299_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0820_  (.Y(\i_ibex/load_store_unit_i/_0300_ ),
    .B1(net1401),
    .B2(data_rdata_i[11]),
    .A2(net1410),
    .A1(data_rdata_i[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0821_  (.Y(\i_ibex/load_store_unit_i/_0301_ ),
    .B1(net1425),
    .B2(data_rdata_i[27]),
    .A2(net1416),
    .A1(data_rdata_i[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0822_  (.A2(\i_ibex/load_store_unit_i/_0301_ ),
    .A1(\i_ibex/load_store_unit_i/_0300_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0302_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(net397),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0824_  (.Y(\i_ibex/load_store_unit_i/_0304_ ),
    .B1(net1425),
    .B2(\i_ibex/load_store_unit_i/rdata_q [19]),
    .A2(net1416),
    .A1(\i_ibex/load_store_unit_i/rdata_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0825_  (.A2(\i_ibex/load_store_unit_i/_0304_ ),
    .A1(\i_ibex/load_store_unit_i/_0300_ ),
    .B1(net1436),
    .X(\i_ibex/load_store_unit_i/_0305_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0826_  (.B(\i_ibex/load_store_unit_i/_0302_ ),
    .C(\i_ibex/load_store_unit_i/_0305_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0827_  (.Y(\i_ibex/load_store_unit_i/_0306_ ),
    .B1(net1402),
    .B2(data_rdata_i[10]),
    .A2(net1413),
    .A1(data_rdata_i[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0828_  (.Y(\i_ibex/load_store_unit_i/_0307_ ),
    .B1(net1430),
    .B2(data_rdata_i[26]),
    .A2(net1420),
    .A1(data_rdata_i[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0829_  (.A2(\i_ibex/load_store_unit_i/_0307_ ),
    .A1(\i_ibex/load_store_unit_i/_0306_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0308_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0830_  (.Y(\i_ibex/load_store_unit_i/_0309_ ),
    .B1(net1430),
    .B2(\i_ibex/load_store_unit_i/rdata_q [18]),
    .A2(net1420),
    .A1(\i_ibex/load_store_unit_i/rdata_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0831_  (.A2(\i_ibex/load_store_unit_i/_0309_ ),
    .A1(\i_ibex/load_store_unit_i/_0306_ ),
    .B1(net1437),
    .X(\i_ibex/load_store_unit_i/_0310_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0832_  (.B(\i_ibex/load_store_unit_i/_0308_ ),
    .C(\i_ibex/load_store_unit_i/_0310_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0833_  (.Y(\i_ibex/load_store_unit_i/_0311_ ),
    .B1(net1400),
    .B2(data_rdata_i[9]),
    .A2(net1409),
    .A1(data_rdata_i[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0834_  (.Y(\i_ibex/load_store_unit_i/_0312_ ),
    .B1(net1423),
    .B2(data_rdata_i[25]),
    .A2(net1415),
    .A1(data_rdata_i[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0835_  (.A2(\i_ibex/load_store_unit_i/_0312_ ),
    .A1(\i_ibex/load_store_unit_i/_0311_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0313_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0836_  (.Y(\i_ibex/load_store_unit_i/_0314_ ),
    .B1(net1423),
    .B2(\i_ibex/load_store_unit_i/rdata_q [17]),
    .A2(net1414),
    .A1(\i_ibex/load_store_unit_i/rdata_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0837_  (.A2(\i_ibex/load_store_unit_i/_0314_ ),
    .A1(\i_ibex/load_store_unit_i/_0311_ ),
    .B1(net1436),
    .X(\i_ibex/load_store_unit_i/_0315_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0838_  (.B(\i_ibex/load_store_unit_i/_0313_ ),
    .C(\i_ibex/load_store_unit_i/_0315_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0839_  (.Y(\i_ibex/load_store_unit_i/_0316_ ),
    .B1(net1402),
    .B2(data_rdata_i[8]),
    .A2(net1412),
    .A1(data_rdata_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0840_  (.Y(\i_ibex/load_store_unit_i/_0317_ ),
    .B1(net1431),
    .B2(data_rdata_i[24]),
    .A2(net1421),
    .A1(data_rdata_i[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0841_  (.A2(\i_ibex/load_store_unit_i/_0317_ ),
    .A1(\i_ibex/load_store_unit_i/_0316_ ),
    .B1(\i_ibex/load_store_unit_i/_0274_ ),
    .X(\i_ibex/load_store_unit_i/_0318_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0842_  (.Y(\i_ibex/load_store_unit_i/_0319_ ),
    .B1(net1431),
    .B2(\i_ibex/load_store_unit_i/rdata_q [16]),
    .A2(net1420),
    .A1(\i_ibex/load_store_unit_i/rdata_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0843_  (.A2(\i_ibex/load_store_unit_i/_0319_ ),
    .A1(\i_ibex/load_store_unit_i/_0316_ ),
    .B1(net1436),
    .X(\i_ibex/load_store_unit_i/_0320_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 \i_ibex/load_store_unit_i/_0844_  (.B(\i_ibex/load_store_unit_i/_0318_ ),
    .C(\i_ibex/load_store_unit_i/_0320_ ),
    .A(net635),
    .Y(\i_ibex/rf_wdata_lsu [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0845_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0321_ ),
    .B(net1458),
    .A(\i_ibex/load_store_unit_i/rdata_offset_q [0]));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0846_  (.Y(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0321_ ),
    .B2(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .A2(net1458),
    .A1(\i_ibex/load_store_unit_i/rdata_offset_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0847_  (.Y(\i_ibex/load_store_unit_i/_0323_ ),
    .B1(net1428),
    .B2(data_rdata_i[23]),
    .A2(net1418),
    .A1(data_rdata_i[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0848_  (.Y(\i_ibex/load_store_unit_i/_0324_ ),
    .A(\i_ibex/load_store_unit_i/_0322_ ),
    .B(\i_ibex/load_store_unit_i/_0323_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0849_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/rdata_q [23]),
    .A2(net1412),
    .Y(\i_ibex/load_store_unit_i/_0325_ ),
    .B1(\i_ibex/load_store_unit_i/_0324_ ));
 sg13g2_or2_1 \i_ibex/load_store_unit_i/_0850_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0326_ ),
    .B(\i_ibex/load_store_unit_i/_0215_ ),
    .A(net1428));
 sg13g2_buf_2 load_slew394 (.A(net891),
    .X(net394),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0852_  (.B1(net1456),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0328_ ),
    .VSS(VSS),
    .A1(data_rdata_i[7]),
    .A2(\i_ibex/load_store_unit_i/_0326_ ));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0853_  (.A(\i_ibex/load_store_unit_i/_0325_ ),
    .B(\i_ibex/load_store_unit_i/_0328_ ),
    .Y(\i_ibex/load_store_unit_i/_0329_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0854_  (.VSS(VSS),
    .VDD(VDD),
    .A1(data_rdata_i[31]),
    .A2(net1412),
    .Y(\i_ibex/load_store_unit_i/_0330_ ),
    .B1(\i_ibex/load_store_unit_i/_0324_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0855_  (.B1(net1457),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0331_ ),
    .VSS(VSS),
    .A1(data_rdata_i[7]),
    .A2(net1399));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0856_  (.A(\i_ibex/load_store_unit_i/_0330_ ),
    .B(\i_ibex/load_store_unit_i/_0331_ ),
    .Y(\i_ibex/load_store_unit_i/_0332_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0857_  (.Y(\i_ibex/load_store_unit_i/_0333_ ),
    .B1(net1430),
    .B2(\i_ibex/load_store_unit_i/rdata_q [15]),
    .A2(net1420),
    .A1(\i_ibex/load_store_unit_i/rdata_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0858_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0334_ ),
    .A(\i_ibex/load_store_unit_i/_0333_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0859_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[7]),
    .C1(\i_ibex/load_store_unit_i/_0334_ ),
    .B1(\i_ibex/load_store_unit_i/_0230_ ),
    .A1(\i_ibex/load_store_unit_i/rdata_q [23]),
    .Y(\i_ibex/load_store_unit_i/_0335_ ),
    .A2(net1412));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0860_  (.A(net1436),
    .B(\i_ibex/load_store_unit_i/_0335_ ),
    .Y(\i_ibex/load_store_unit_i/_0336_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_2 \i_ibex/load_store_unit_i/_0861_  (.A(\i_ibex/load_store_unit_i/_0329_ ),
    .B(\i_ibex/load_store_unit_i/_0332_ ),
    .C(\i_ibex/load_store_unit_i/_0336_ ),
    .X(\i_ibex/rf_wdata_lsu [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0862_  (.Y(\i_ibex/load_store_unit_i/_0337_ ),
    .B1(net1423),
    .B2(\i_ibex/load_store_unit_i/rdata_q [14]),
    .A2(net1414),
    .A1(\i_ibex/load_store_unit_i/rdata_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0863_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0338_ ),
    .A(\i_ibex/load_store_unit_i/_0337_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0864_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[6]),
    .C1(\i_ibex/load_store_unit_i/_0338_ ),
    .B1(net1400),
    .A1(\i_ibex/load_store_unit_i/rdata_q [22]),
    .Y(\i_ibex/load_store_unit_i/_0339_ ),
    .A2(net1409));
 sg13g2_or2_2 \i_ibex/load_store_unit_i/_0865_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/load_store_unit_i/_0340_ ),
    .B(net1458),
    .A(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ));
 sg13g2_buf_2 fanout393 (.A(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .X(net393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0867_  (.Y(\i_ibex/load_store_unit_i/_0342_ ),
    .B1(net1456),
    .B2(\i_ibex/load_store_unit_i/rdata_q [22]),
    .A2(net1457),
    .A1(data_rdata_i[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0868_  (.Y(\i_ibex/load_store_unit_i/_0343_ ),
    .B1(net1424),
    .B2(data_rdata_i[22]),
    .A2(net1415),
    .A1(data_rdata_i[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 \i_ibex/load_store_unit_i/_0869_  (.A(net1457),
    .B(net1456),
    .Y(\i_ibex/load_store_unit_i/_0344_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0870_  (.A2(\i_ibex/load_store_unit_i/_0343_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0345_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0871_  (.B1(\i_ibex/load_store_unit_i/_0345_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0346_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0342_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0872_  (.B1(\i_ibex/load_store_unit_i/_0346_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0347_ ),
    .VSS(VSS),
    .A1(data_rdata_i[6]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0873_  (.B1(\i_ibex/load_store_unit_i/_0347_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [6]),
    .VSS(VSS),
    .A1(net1435),
    .A2(\i_ibex/load_store_unit_i/_0339_ ));
 sg13g2_buf_2 fanout392 (.A(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .X(net392),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout391 (.A(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .X(net391),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0876_  (.Y(\i_ibex/load_store_unit_i/_0350_ ),
    .B1(net1426),
    .B2(\i_ibex/load_store_unit_i/rdata_q [13]),
    .A2(net1417),
    .A1(\i_ibex/load_store_unit_i/rdata_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0877_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0351_ ),
    .A(\i_ibex/load_store_unit_i/_0350_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0878_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[5]),
    .C1(\i_ibex/load_store_unit_i/_0351_ ),
    .B1(\i_ibex/load_store_unit_i/_0216_ ),
    .A1(\i_ibex/load_store_unit_i/rdata_q [21]),
    .Y(\i_ibex/load_store_unit_i/_0352_ ),
    .A2(net1410));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0879_  (.Y(\i_ibex/load_store_unit_i/_0353_ ),
    .B1(net1456),
    .B2(\i_ibex/load_store_unit_i/rdata_q [21]),
    .A2(net1457),
    .A1(data_rdata_i[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0880_  (.Y(\i_ibex/load_store_unit_i/_0354_ ),
    .B1(net1425),
    .B2(data_rdata_i[21]),
    .A2(net1416),
    .A1(data_rdata_i[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0881_  (.A2(\i_ibex/load_store_unit_i/_0354_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0355_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0882_  (.B1(\i_ibex/load_store_unit_i/_0355_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0356_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0353_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0883_  (.B1(\i_ibex/load_store_unit_i/_0356_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0357_ ),
    .VSS(VSS),
    .A1(data_rdata_i[5]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0884_  (.B1(\i_ibex/load_store_unit_i/_0357_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [5]),
    .VSS(VSS),
    .A1(net1436),
    .A2(\i_ibex/load_store_unit_i/_0352_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0885_  (.Y(\i_ibex/load_store_unit_i/_0358_ ),
    .B1(net1424),
    .B2(\i_ibex/load_store_unit_i/rdata_q [12]),
    .A2(net1415),
    .A1(\i_ibex/load_store_unit_i/rdata_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0886_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0359_ ),
    .A(\i_ibex/load_store_unit_i/_0358_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0887_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[4]),
    .C1(\i_ibex/load_store_unit_i/_0359_ ),
    .B1(net1401),
    .A1(\i_ibex/load_store_unit_i/rdata_q [20]),
    .Y(\i_ibex/load_store_unit_i/_0360_ ),
    .A2(net1409));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0888_  (.Y(\i_ibex/load_store_unit_i/_0361_ ),
    .B1(net1456),
    .B2(\i_ibex/load_store_unit_i/rdata_q [20]),
    .A2(net1457),
    .A1(data_rdata_i[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0889_  (.Y(\i_ibex/load_store_unit_i/_0362_ ),
    .B1(net1424),
    .B2(data_rdata_i[20]),
    .A2(net1415),
    .A1(data_rdata_i[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0890_  (.A2(\i_ibex/load_store_unit_i/_0362_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0363_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0891_  (.B1(\i_ibex/load_store_unit_i/_0363_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0364_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0361_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0892_  (.B1(\i_ibex/load_store_unit_i/_0364_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0365_ ),
    .VSS(VSS),
    .A1(data_rdata_i[4]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0893_  (.B1(\i_ibex/load_store_unit_i/_0365_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [4]),
    .VSS(VSS),
    .A1(net1435),
    .A2(\i_ibex/load_store_unit_i/_0360_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0894_  (.Y(\i_ibex/load_store_unit_i/_0366_ ),
    .B1(net1425),
    .B2(\i_ibex/load_store_unit_i/rdata_q [11]),
    .A2(net1416),
    .A1(\i_ibex/load_store_unit_i/rdata_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0895_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0367_ ),
    .A(\i_ibex/load_store_unit_i/_0366_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0896_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[3]),
    .C1(\i_ibex/load_store_unit_i/_0367_ ),
    .B1(net1401),
    .A1(\i_ibex/load_store_unit_i/rdata_q [19]),
    .Y(\i_ibex/load_store_unit_i/_0368_ ),
    .A2(net1410));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0897_  (.Y(\i_ibex/load_store_unit_i/_0369_ ),
    .B1(net1456),
    .B2(\i_ibex/load_store_unit_i/rdata_q [19]),
    .A2(net1457),
    .A1(data_rdata_i[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0898_  (.Y(\i_ibex/load_store_unit_i/_0370_ ),
    .B1(net1425),
    .B2(data_rdata_i[19]),
    .A2(net1416),
    .A1(data_rdata_i[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0899_  (.A2(\i_ibex/load_store_unit_i/_0370_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0371_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0900_  (.B1(\i_ibex/load_store_unit_i/_0371_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0372_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0369_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0901_  (.B1(\i_ibex/load_store_unit_i/_0372_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0373_ ),
    .VSS(VSS),
    .A1(data_rdata_i[3]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0902_  (.B1(\i_ibex/load_store_unit_i/_0373_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [3]),
    .VSS(VSS),
    .A1(net1436),
    .A2(\i_ibex/load_store_unit_i/_0368_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0903_  (.Y(\i_ibex/load_store_unit_i/_0374_ ),
    .B1(net1430),
    .B2(\i_ibex/load_store_unit_i/rdata_q [10]),
    .A2(net1420),
    .A1(\i_ibex/load_store_unit_i/rdata_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0904_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0375_ ),
    .A(\i_ibex/load_store_unit_i/_0374_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0905_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[2]),
    .C1(\i_ibex/load_store_unit_i/_0375_ ),
    .B1(net1402),
    .A1(\i_ibex/load_store_unit_i/rdata_q [18]),
    .Y(\i_ibex/load_store_unit_i/_0376_ ),
    .A2(net1413));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0906_  (.Y(\i_ibex/load_store_unit_i/_0377_ ),
    .B1(\i_ibex/load_store_unit_i/_0242_ ),
    .B2(\i_ibex/load_store_unit_i/rdata_q [18]),
    .A2(\i_ibex/load_store_unit_i/_0235_ ),
    .A1(data_rdata_i[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0907_  (.Y(\i_ibex/load_store_unit_i/_0378_ ),
    .B1(net1424),
    .B2(data_rdata_i[18]),
    .A2(net1415),
    .A1(data_rdata_i[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0908_  (.A2(\i_ibex/load_store_unit_i/_0378_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0379_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0909_  (.B1(\i_ibex/load_store_unit_i/_0379_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0380_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0377_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0910_  (.B1(\i_ibex/load_store_unit_i/_0380_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0381_ ),
    .VSS(VSS),
    .A1(data_rdata_i[2]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0911_  (.B1(\i_ibex/load_store_unit_i/_0381_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [2]),
    .VSS(VSS),
    .A1(net1437),
    .A2(\i_ibex/load_store_unit_i/_0376_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0912_  (.Y(\i_ibex/load_store_unit_i/_0382_ ),
    .B1(net1411),
    .B2(data_rdata_i[20]),
    .A2(net1428),
    .A1(data_rdata_i[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0913_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0383_ ),
    .A(\i_ibex/load_store_unit_i/_0382_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0914_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[28]),
    .C1(\i_ibex/load_store_unit_i/_0383_ ),
    .B1(net1403),
    .A1(data_rdata_i[4]),
    .Y(\i_ibex/load_store_unit_i/_0384_ ),
    .A2(net1418));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0915_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [28]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0384_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0916_  (.Y(\i_ibex/load_store_unit_i/_0385_ ),
    .B1(net1425),
    .B2(\i_ibex/load_store_unit_i/rdata_q [9]),
    .A2(net1416),
    .A1(\i_ibex/load_store_unit_i/rdata_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0917_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0386_ ),
    .A(\i_ibex/load_store_unit_i/_0385_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0918_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[1]),
    .C1(\i_ibex/load_store_unit_i/_0386_ ),
    .B1(net1401),
    .A1(\i_ibex/load_store_unit_i/rdata_q [17]),
    .Y(\i_ibex/load_store_unit_i/_0387_ ),
    .A2(net1410));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0919_  (.Y(\i_ibex/load_store_unit_i/_0388_ ),
    .B1(net1456),
    .B2(\i_ibex/load_store_unit_i/rdata_q [17]),
    .A2(net1457),
    .A1(data_rdata_i[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0920_  (.Y(\i_ibex/load_store_unit_i/_0389_ ),
    .B1(net1424),
    .B2(data_rdata_i[17]),
    .A2(net1415),
    .A1(data_rdata_i[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0921_  (.A2(\i_ibex/load_store_unit_i/_0389_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0390_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0922_  (.B1(\i_ibex/load_store_unit_i/_0390_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0391_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0388_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0923_  (.B1(\i_ibex/load_store_unit_i/_0391_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0392_ ),
    .VSS(VSS),
    .A1(data_rdata_i[1]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0924_  (.B1(\i_ibex/load_store_unit_i/_0392_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [1]),
    .VSS(VSS),
    .A1(net1436),
    .A2(\i_ibex/load_store_unit_i/_0387_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0925_  (.Y(\i_ibex/load_store_unit_i/_0393_ ),
    .B1(net1431),
    .B2(\i_ibex/load_store_unit_i/rdata_q [8]),
    .A2(net1421),
    .A1(\i_ibex/load_store_unit_i/rdata_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0926_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0394_ ),
    .A(\i_ibex/load_store_unit_i/_0393_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0927_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[0]),
    .C1(\i_ibex/load_store_unit_i/_0394_ ),
    .B1(net1403),
    .A1(\i_ibex/load_store_unit_i/rdata_q [16]),
    .Y(\i_ibex/load_store_unit_i/_0395_ ),
    .A2(net1413));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0928_  (.Y(\i_ibex/load_store_unit_i/_0396_ ),
    .B1(\i_ibex/load_store_unit_i/_0242_ ),
    .B2(\i_ibex/load_store_unit_i/rdata_q [16]),
    .A2(\i_ibex/load_store_unit_i/_0235_ ),
    .A1(data_rdata_i[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0929_  (.Y(\i_ibex/load_store_unit_i/_0397_ ),
    .B1(net1430),
    .B2(data_rdata_i[16]),
    .A2(net1420),
    .A1(data_rdata_i[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 \i_ibex/load_store_unit_i/_0930_  (.A2(\i_ibex/load_store_unit_i/_0397_ ),
    .A1(\i_ibex/load_store_unit_i/_0322_ ),
    .B1(\i_ibex/load_store_unit_i/_0344_ ),
    .X(\i_ibex/load_store_unit_i/_0398_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0931_  (.B1(\i_ibex/load_store_unit_i/_0398_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0399_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0340_ ),
    .A2(\i_ibex/load_store_unit_i/_0396_ ));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0932_  (.B1(\i_ibex/load_store_unit_i/_0399_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0400_ ),
    .VSS(VSS),
    .A1(data_rdata_i[0]),
    .A2(net1399));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0933_  (.B1(\i_ibex/load_store_unit_i/_0400_ ),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [0]),
    .VSS(VSS),
    .A1(net1437),
    .A2(\i_ibex/load_store_unit_i/_0395_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0934_  (.Y(\i_ibex/load_store_unit_i/_0401_ ),
    .B1(net1410),
    .B2(data_rdata_i[19]),
    .A2(net1425),
    .A1(data_rdata_i[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0935_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0402_ ),
    .A(\i_ibex/load_store_unit_i/_0401_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0936_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[27]),
    .C1(\i_ibex/load_store_unit_i/_0402_ ),
    .B1(net1401),
    .A1(data_rdata_i[3]),
    .Y(\i_ibex/load_store_unit_i/_0403_ ),
    .A2(net1416));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0937_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [27]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0403_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0938_  (.Y(\i_ibex/load_store_unit_i/_0404_ ),
    .B1(net1413),
    .B2(data_rdata_i[18]),
    .A2(net1428),
    .A1(data_rdata_i[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0939_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0405_ ),
    .A(\i_ibex/load_store_unit_i/_0404_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0940_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[26]),
    .C1(\i_ibex/load_store_unit_i/_0405_ ),
    .B1(net1402),
    .A1(data_rdata_i[2]),
    .Y(\i_ibex/load_store_unit_i/_0406_ ),
    .A2(net1418));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0941_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [26]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0406_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0942_  (.Y(\i_ibex/load_store_unit_i/_0407_ ),
    .B1(net1409),
    .B2(data_rdata_i[17]),
    .A2(net1423),
    .A1(data_rdata_i[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0943_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0408_ ),
    .A(\i_ibex/load_store_unit_i/_0407_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0944_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[25]),
    .C1(\i_ibex/load_store_unit_i/_0408_ ),
    .B1(net1400),
    .A1(data_rdata_i[1]),
    .Y(\i_ibex/load_store_unit_i/_0409_ ),
    .A2(net1414));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0945_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [25]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0409_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0946_  (.Y(\i_ibex/load_store_unit_i/_0410_ ),
    .B1(net1413),
    .B2(data_rdata_i[16]),
    .A2(net1430),
    .A1(data_rdata_i[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0947_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0411_ ),
    .A(\i_ibex/load_store_unit_i/_0410_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0948_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[24]),
    .C1(\i_ibex/load_store_unit_i/_0411_ ),
    .B1(net1402),
    .A1(data_rdata_i[0]),
    .Y(\i_ibex/load_store_unit_i/_0412_ ),
    .A2(net1420));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0949_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [24]),
    .VSS(VSS),
    .A1(net1433),
    .A2(\i_ibex/load_store_unit_i/_0412_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0950_  (.Y(\i_ibex/load_store_unit_i/_0413_ ),
    .B1(net1429),
    .B2(data_rdata_i[7]),
    .A2(net1419),
    .A1(\i_ibex/load_store_unit_i/rdata_q [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0951_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0414_ ),
    .A(\i_ibex/load_store_unit_i/_0413_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0952_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[23]),
    .C1(\i_ibex/load_store_unit_i/_0414_ ),
    .B1(net1403),
    .A1(data_rdata_i[15]),
    .Y(\i_ibex/load_store_unit_i/_0415_ ),
    .A2(net1412));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0953_  (.B1(net1276),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [23]),
    .VSS(VSS),
    .A1(net1434),
    .A2(\i_ibex/load_store_unit_i/_0415_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0954_  (.Y(\i_ibex/load_store_unit_i/_0416_ ),
    .B1(net1409),
    .B2(data_rdata_i[14]),
    .A2(net1414),
    .A1(\i_ibex/load_store_unit_i/rdata_q [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/load_store_unit_i/_0955_  (.VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0417_ ),
    .A(\i_ibex/load_store_unit_i/_0416_ ),
    .VSS(VSS));
 sg13g2_a221oi_1 \i_ibex/load_store_unit_i/_0956_  (.VSS(VSS),
    .VDD(VDD),
    .B2(data_rdata_i[22]),
    .C1(\i_ibex/load_store_unit_i/_0417_ ),
    .B1(net1400),
    .A1(data_rdata_i[6]),
    .Y(\i_ibex/load_store_unit_i/_0418_ ),
    .A2(net1423));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0957_  (.B1(net1277),
    .VDD(VDD),
    .Y(\i_ibex/rf_wdata_lsu [22]),
    .VSS(VSS),
    .A1(net1432),
    .A2(\i_ibex/load_store_unit_i/_0418_ ));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0958_  (.Y(\i_ibex/load_store_unit_i/_0419_ ),
    .B(data_rvalid_i),
    .A_N(data_err_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 \i_ibex/load_store_unit_i/_0959_  (.A(\i_ibex/load_store_unit_i/pmp_err_q ),
    .B(\i_ibex/load_store_unit_i/lsu_err_q ),
    .C(\i_ibex/load_store_unit_i/_0419_ ),
    .D(\i_ibex/load_store_unit_i/_0182_ ),
    .Y(\i_ibex/rf_we_lsu ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0960_  (.A(\i_ibex/lsu_we ),
    .B(\i_ibex/load_store_unit_i/_0123_ ),
    .Y(\i_ibex/perf_load ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 \i_ibex/load_store_unit_i/_0961_  (.X(\i_ibex/perf_store ),
    .A(\i_ibex/lsu_req ),
    .B(\i_ibex/lsu_we ),
    .C(\i_ibex/load_store_unit_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 \i_ibex/load_store_unit_i/_0962_  (.A(net1460),
    .B_N(\i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ),
    .Y(\i_ibex/load_store_unit_i/_0420_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0963_  (.B1(\i_ibex/load_store_unit_i/_0091_ ),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0421_ ),
    .VSS(VSS),
    .A1(\i_ibex/load_store_unit_i/_0201_ ),
    .A2(\i_ibex/load_store_unit_i/_0420_ ));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0964_  (.Y(\i_ibex/load_store_unit_i/_0422_ ),
    .A(net1769),
    .B(\i_ibex/load_store_unit_i/_0072_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0965_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/_0421_ ),
    .A2(\i_ibex/load_store_unit_i/_0422_ ),
    .Y(\i_ibex/load_store_unit_i/_0423_ ),
    .B1(net1462));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0966_  (.Y(\i_ibex/load_store_unit_i/_0424_ ),
    .B(\i_ibex/load_store_unit_i/_0423_ ),
    .A_N(\i_ibex/load_store_unit_i/_0190_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 \i_ibex/load_store_unit_i/_0967_  (.Y(\i_ibex/load_store_unit_i/_0425_ ),
    .B(\i_ibex/load_store_unit_i/_0092_ ),
    .A_N(\i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0968_  (.Y(\i_ibex/load_store_unit_i/_0426_ ),
    .A(\i_ibex/load_store_unit_i/_0425_ ),
    .B(\i_ibex/load_store_unit_i/_0189_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 \i_ibex/load_store_unit_i/_0969_  (.B1(net45),
    .VDD(VDD),
    .Y(\i_ibex/load_store_unit_i/_0427_ ),
    .VSS(VSS),
    .A1(\i_ibex/lsu_req ),
    .A2(\i_ibex/load_store_unit_i/_0426_ ));
 sg13g2_a22oi_1 \i_ibex/load_store_unit_i/_0970_  (.Y(\i_ibex/load_store_unit_i/_0041_ ),
    .B1(\i_ibex/load_store_unit_i/_0427_ ),
    .B2(\i_ibex/load_store_unit_i/_0423_ ),
    .A2(\i_ibex/load_store_unit_i/_0424_ ),
    .A1(\i_ibex/load_store_unit_i/_0080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0971_  (.A0(\i_ibex/load_store_unit_i/rdata_offset_q [0]),
    .A1(net472),
    .S(\i_ibex/load_store_unit_i/_0129_ ),
    .X(\i_ibex/load_store_unit_i/_0042_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0972_  (.A0(\i_ibex/load_store_unit_i/rdata_offset_q [1]),
    .A1(net434),
    .S(\i_ibex/load_store_unit_i/_0129_ ),
    .X(\i_ibex/load_store_unit_i/_0043_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 \i_ibex/load_store_unit_i/_0973_  (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_ibex/load_store_unit_i/pmp_err_q ),
    .A2(\i_ibex/load_store_unit_i/_0425_ ),
    .Y(\i_ibex/load_store_unit_i/_0428_ ),
    .B1(net1785));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_0974_  (.Y(\i_ibex/load_store_unit_i/_0429_ ),
    .A(\i_ibex/load_store_unit_i/lsu_rdata_valid_o_$_AND__Y_B ),
    .B(\i_ibex/load_store_unit_i/_0426_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 \i_ibex/load_store_unit_i/_0975_  (.A(\i_ibex/load_store_unit_i/_0428_ ),
    .B(\i_ibex/load_store_unit_i/_0429_ ),
    .Y(\i_ibex/load_store_unit_i/_0430_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout390 (.A(\i_ibex/cs_registers_i/mhpmcounterh_we [2]),
    .X(net390),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0977_  (.A0(\i_ibex/load_store_unit_i/rdata_q [0]),
    .A1(net1706),
    .S(net1319),
    .X(\i_ibex/load_store_unit_i/_0044_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0978_  (.A0(\i_ibex/load_store_unit_i/rdata_q [10]),
    .A1(net1731),
    .S(net1319),
    .X(\i_ibex/load_store_unit_i/_0045_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0979_  (.A0(\i_ibex/load_store_unit_i/rdata_q [11]),
    .A1(net1727),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0046_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0980_  (.A0(\i_ibex/load_store_unit_i/rdata_q [12]),
    .A1(net1704),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0047_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0981_  (.A0(\i_ibex/load_store_unit_i/rdata_q [13]),
    .A1(net1717),
    .S(net1319),
    .X(\i_ibex/load_store_unit_i/_0048_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0982_  (.A0(\i_ibex/load_store_unit_i/rdata_q [14]),
    .A1(net1711),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0983_  (.A0(\i_ibex/load_store_unit_i/rdata_q [15]),
    .A1(net1750),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0050_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0984_  (.A0(\i_ibex/load_store_unit_i/rdata_q [16]),
    .A1(net1741),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0051_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0985_  (.A0(\i_ibex/load_store_unit_i/rdata_q [17]),
    .A1(net1725),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0986_  (.A0(\i_ibex/load_store_unit_i/rdata_q [18]),
    .A1(net1745),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0053_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout389 (.X(net389),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0226_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0988_  (.A0(\i_ibex/load_store_unit_i/rdata_q [19]),
    .A1(net1720),
    .S(net1317),
    .X(\i_ibex/load_store_unit_i/_0054_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0989_  (.A0(\i_ibex/load_store_unit_i/rdata_q [1]),
    .A1(net1746),
    .S(net1317),
    .X(\i_ibex/load_store_unit_i/_0055_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0990_  (.A0(\i_ibex/load_store_unit_i/rdata_q [20]),
    .A1(net1694),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0056_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0991_  (.A0(\i_ibex/load_store_unit_i/rdata_q [21]),
    .A1(net1729),
    .S(net1319),
    .X(\i_ibex/load_store_unit_i/_0057_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0992_  (.A0(\i_ibex/load_store_unit_i/rdata_q [22]),
    .A1(net1739),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0058_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0993_  (.A0(\i_ibex/load_store_unit_i/rdata_q [23]),
    .A1(net1744),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0059_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0994_  (.A0(\i_ibex/load_store_unit_i/rdata_q [2]),
    .A1(net1736),
    .S(net1317),
    .X(\i_ibex/load_store_unit_i/_0060_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0995_  (.A0(\i_ibex/load_store_unit_i/rdata_q [3]),
    .A1(net1733),
    .S(net1317),
    .X(\i_ibex/load_store_unit_i/_0061_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0996_  (.A0(\i_ibex/load_store_unit_i/rdata_q [4]),
    .A1(net1742),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0062_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0997_  (.A0(\i_ibex/load_store_unit_i/rdata_q [5]),
    .A1(net1713),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0063_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0998_  (.A0(\i_ibex/load_store_unit_i/rdata_q [6]),
    .A1(net1715),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0064_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_0999_  (.A0(\i_ibex/load_store_unit_i/rdata_q [7]),
    .A1(net1752),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0065_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_1000_  (.A0(\i_ibex/load_store_unit_i/rdata_q [8]),
    .A1(net1748),
    .S(net1318),
    .X(\i_ibex/load_store_unit_i/_0066_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 \i_ibex/load_store_unit_i/_1001_  (.A0(\i_ibex/load_store_unit_i/rdata_q [9]),
    .A1(net1722),
    .S(net1316),
    .X(\i_ibex/load_store_unit_i/_0067_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 \i_ibex/load_store_unit_i/_1002_  (.Y(\i_ibex/load_store_unit_i/_0433_ ),
    .A(\i_ibex/load_store_unit_i/data_we_q ),
    .B(\i_ibex/load_store_unit_i/_0105_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 \i_ibex/load_store_unit_i/_1003_  (.VSS(VSS),
    .VDD(VDD),
    .B1(\i_ibex/load_store_unit_i/_0433_ ),
    .Y(\i_ibex/lsu_store_err ),
    .A2(\i_ibex/load_store_unit_i/_0181_ ),
    .A1(\i_ibex/load_store_unit_i/_0080_ ));
 sg13g2_tiehi \i_ibex/cs_registers_i/u_mtvec_csr/_073__381  (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net381));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0000_ ),
    .Q(\i_ibex/lsu_addr_last [0]),
    .Q_N(\i_ibex/load_store_unit_i/_0491_ ),
    .CLK(clknet_leaf_106_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[10]_reg  (.CLK(clknet_leaf_97_clk_i_regs),
    .RESET_B(net1565),
    .D(\i_ibex/load_store_unit_i/_0001_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0490_ ),
    .Q(\i_ibex/lsu_addr_last [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[11]_reg  (.CLK(clknet_leaf_97_clk_i_regs),
    .RESET_B(net1564),
    .D(\i_ibex/load_store_unit_i/_0002_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0489_ ),
    .Q(\i_ibex/lsu_addr_last [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[12]_reg  (.CLK(clknet_leaf_96_clk_i_regs),
    .RESET_B(net1565),
    .D(\i_ibex/load_store_unit_i/_0003_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0488_ ),
    .Q(\i_ibex/lsu_addr_last [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[13]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1564),
    .D(\i_ibex/load_store_unit_i/_0004_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0487_ ),
    .Q(\i_ibex/lsu_addr_last [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[14]_reg  (.CLK(clknet_leaf_97_clk_i_regs),
    .RESET_B(net1564),
    .D(\i_ibex/load_store_unit_i/_0005_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0486_ ),
    .Q(\i_ibex/lsu_addr_last [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[15]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1563),
    .D(\i_ibex/load_store_unit_i/_0006_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0485_ ),
    .Q(\i_ibex/lsu_addr_last [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[16]_reg  (.RESET_B(net1565),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0007_ ),
    .Q(\i_ibex/lsu_addr_last [16]),
    .Q_N(\i_ibex/load_store_unit_i/_0484_ ),
    .CLK(clknet_leaf_96_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[17]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1563),
    .D(\i_ibex/load_store_unit_i/_0008_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0483_ ),
    .Q(\i_ibex/lsu_addr_last [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[18]_reg  (.RESET_B(net1566),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0009_ ),
    .Q(\i_ibex/lsu_addr_last [18]),
    .Q_N(\i_ibex/load_store_unit_i/_0482_ ),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[19]_reg  (.RESET_B(net1565),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0010_ ),
    .Q(\i_ibex/lsu_addr_last [19]),
    .Q_N(\i_ibex/load_store_unit_i/_0481_ ),
    .CLK(clknet_leaf_96_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[1]_reg  (.RESET_B(net1664),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0011_ ),
    .Q(\i_ibex/lsu_addr_last [1]),
    .Q_N(\i_ibex/load_store_unit_i/_0480_ ),
    .CLK(clknet_leaf_106_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[20]_reg  (.RESET_B(net1563),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0012_ ),
    .Q(\i_ibex/lsu_addr_last [20]),
    .Q_N(\i_ibex/load_store_unit_i/_0479_ ),
    .CLK(clknet_leaf_99_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[21]_reg  (.RESET_B(net1566),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0013_ ),
    .Q(\i_ibex/lsu_addr_last [21]),
    .Q_N(\i_ibex/load_store_unit_i/_0478_ ),
    .CLK(clknet_leaf_99_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[22]_reg  (.CLK(clknet_leaf_99_clk_i_regs),
    .RESET_B(net1563),
    .D(\i_ibex/load_store_unit_i/_0014_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0477_ ),
    .Q(\i_ibex/lsu_addr_last [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[23]_reg  (.CLK(clknet_5_16__leaf_clk_i_regs),
    .RESET_B(net1566),
    .D(\i_ibex/load_store_unit_i/_0015_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0476_ ),
    .Q(\i_ibex/lsu_addr_last [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[24]_reg  (.RESET_B(net1566),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0016_ ),
    .Q(\i_ibex/lsu_addr_last [24]),
    .Q_N(\i_ibex/load_store_unit_i/_0475_ ),
    .CLK(clknet_leaf_99_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[25]_reg  (.CLK(clknet_leaf_99_clk_i_regs),
    .RESET_B(net1563),
    .D(\i_ibex/load_store_unit_i/_0017_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0474_ ),
    .Q(\i_ibex/lsu_addr_last [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[26]_reg  (.CLK(clknet_leaf_36_clk_i_regs),
    .RESET_B(net1566),
    .D(\i_ibex/load_store_unit_i/_0018_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0473_ ),
    .Q(\i_ibex/lsu_addr_last [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[27]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1563),
    .D(\i_ibex/load_store_unit_i/_0019_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0472_ ),
    .Q(\i_ibex/lsu_addr_last [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[28]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1564),
    .D(\i_ibex/load_store_unit_i/_0020_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0471_ ),
    .Q(\i_ibex/lsu_addr_last [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[29]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1564),
    .D(\i_ibex/load_store_unit_i/_0021_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0470_ ),
    .Q(\i_ibex/lsu_addr_last [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[2]_reg  (.CLK(clknet_5_29__leaf_clk_i_regs),
    .RESET_B(net1576),
    .D(\i_ibex/load_store_unit_i/_0022_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0469_ ),
    .Q(\i_ibex/lsu_addr_last [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/addr_last_o[30]_reg  (.RESET_B(net1563),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0023_ ),
    .Q(\i_ibex/lsu_addr_last [30]),
    .Q_N(\i_ibex/load_store_unit_i/_0468_ ),
    .CLK(clknet_leaf_99_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[31]_reg  (.CLK(clknet_leaf_99_clk_i_regs),
    .RESET_B(net1563),
    .D(\i_ibex/load_store_unit_i/_0024_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0467_ ),
    .Q(\i_ibex/lsu_addr_last [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[3]_reg  (.CLK(clknet_leaf_83_clk_i_regs),
    .RESET_B(net1575),
    .D(\i_ibex/load_store_unit_i/_0025_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0466_ ),
    .Q(\i_ibex/lsu_addr_last [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[4]_reg  (.CLK(clknet_leaf_92_clk_i_regs),
    .RESET_B(net1578),
    .D(\i_ibex/load_store_unit_i/_0026_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0465_ ),
    .Q(\i_ibex/lsu_addr_last [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[5]_reg  (.CLK(clknet_leaf_92_clk_i_regs),
    .RESET_B(net1575),
    .D(\i_ibex/load_store_unit_i/_0027_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0464_ ),
    .Q(\i_ibex/lsu_addr_last [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[6]_reg  (.CLK(clknet_leaf_91_clk_i_regs),
    .RESET_B(net1578),
    .D(\i_ibex/load_store_unit_i/_0028_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0463_ ),
    .Q(\i_ibex/lsu_addr_last [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[7]_reg  (.CLK(clknet_leaf_93_clk_i_regs),
    .RESET_B(net1575),
    .D(\i_ibex/load_store_unit_i/_0029_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0462_ ),
    .Q(\i_ibex/lsu_addr_last [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[8]_reg  (.CLK(clknet_leaf_91_clk_i_regs),
    .RESET_B(net1575),
    .D(\i_ibex/load_store_unit_i/_0030_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0461_ ),
    .Q(\i_ibex/lsu_addr_last [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/addr_last_o[9]_reg  (.CLK(clknet_leaf_98_clk_i_regs),
    .RESET_B(net1564),
    .D(\i_ibex/load_store_unit_i/_0031_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0460_ ),
    .Q(\i_ibex/lsu_addr_last [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/data_sign_ext_q_reg  (.CLK(clknet_leaf_135_clk_i_regs),
    .RESET_B(net1657),
    .D(\i_ibex/load_store_unit_i/_0032_ ),
    .Q_N(\i_ibex/load_store_unit_i/_0459_ ),
    .Q(\i_ibex/load_store_unit_i/data_sign_ext_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/data_type_q[0]_reg  (.CLK(clknet_leaf_135_clk_i_regs),
    .RESET_B(net1657),
    .D(\i_ibex/load_store_unit_i/_0033_ ),
    .Q_N(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_Y ),
    .Q(\i_ibex/load_store_unit_i/data_type_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/data_type_q[1]_reg  (.CLK(clknet_leaf_135_clk_i_regs),
    .RESET_B(net1657),
    .D(\i_ibex/load_store_unit_i/_0034_ ),
    .Q_N(\i_ibex/load_store_unit_i/data_type_q_$_NOT__A_1_Y ),
    .Q(\i_ibex/load_store_unit_i/data_type_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/data_we_q_reg  (.CLK(clknet_leaf_104_clk_i_regs),
    .RESET_B(rst_ni),
    .D(\i_ibex/load_store_unit_i/_0035_ ),
    .Q_N(\i_ibex/load_store_unit_i/lsu_rdata_valid_o_$_AND__Y_B ),
    .Q(\i_ibex/load_store_unit_i/data_we_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/handle_misaligned_q_reg  (.CLK(clknet_leaf_105_clk_i_regs),
    .RESET_B(net1664),
    .D(\i_ibex/load_store_unit_i/_0036_ ),
    .Q_N(\i_ibex/load_store_unit_i/data_be_o_$_MUX__Y_A [3]),
    .Q(\i_ibex/load_store_unit_i/handle_misaligned_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg  (.CLK(clknet_leaf_103_clk_i_regs),
    .RESET_B(net1657),
    .D(net1756),
    .Q_N(\i_ibex/load_store_unit_i/ls_fsm_cs[0]_reg_E_$_AND__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .Q(\i_ibex/load_store_unit_i/ls_fsm_cs [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/ls_fsm_cs[1]_reg  (.RESET_B(net1657),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0038_ ),
    .Q(\i_ibex/load_store_unit_i/ls_fsm_cs [1]),
    .Q_N(\i_ibex/load_store_unit_i/busy_o_$_NOT__A_Y_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_103_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/ls_fsm_cs[2]_reg  (.RESET_B(net1657),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0039_ ),
    .Q(\i_ibex/load_store_unit_i/ls_fsm_cs [2]),
    .Q_N(\i_ibex/load_store_unit_i/busy_o_$_OR__Y_A_$_OR__A_B ),
    .CLK(clknet_leaf_104_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/lsu_err_q_reg  (.CLK(clknet_leaf_103_clk_i_regs),
    .RESET_B(net1664),
    .D(net1758),
    .Q_N(\i_ibex/load_store_unit_i/lsu_err_q_$_NOT__A_Y ),
    .Q(\i_ibex/load_store_unit_i/lsu_err_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/pmp_err_q_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0041_ ),
    .Q(\i_ibex/load_store_unit_i/pmp_err_q ),
    .Q_N(\i_ibex/load_store_unit_i/_0458_ ),
    .CLK(clknet_leaf_113_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_offset_q[0]_reg  (.RESET_B(net1657),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0042_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_offset_q [0]),
    .Q_N(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_Y ),
    .CLK(clknet_5_16__leaf_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_offset_q[1]_reg  (.CLK(clknet_leaf_135_clk_i_regs),
    .RESET_B(net1657),
    .D(\i_ibex/load_store_unit_i/_0043_ ),
    .Q_N(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_1_Y ),
    .Q(\i_ibex/load_store_unit_i/rdata_offset_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[0]_reg  (.CLK(clknet_leaf_130_clk_i_regs),
    .RESET_B(net1658),
    .D(net1707),
    .Q_N(\i_ibex/load_store_unit_i/_0457_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[10]_reg  (.CLK(clknet_leaf_130_clk_i_regs),
    .RESET_B(net1658),
    .D(net1732),
    .Q_N(\i_ibex/load_store_unit_i/_0456_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[11]_reg  (.CLK(clknet_leaf_132_clk_i_regs),
    .RESET_B(net1580),
    .D(net1728),
    .Q_N(\i_ibex/load_store_unit_i/_0455_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[12]_reg  (.CLK(clknet_leaf_134_clk_i_regs),
    .RESET_B(net1659),
    .D(net1705),
    .Q_N(\i_ibex/load_store_unit_i/_0454_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[13]_reg  (.CLK(clknet_leaf_130_clk_i_regs),
    .RESET_B(net1659),
    .D(net1718),
    .Q_N(\i_ibex/load_store_unit_i/_0453_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[14]_reg  (.CLK(clknet_leaf_133_clk_i_regs),
    .RESET_B(net1580),
    .D(net1712),
    .Q_N(\i_ibex/load_store_unit_i/_0452_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[15]_reg  (.CLK(clknet_leaf_135_clk_i_regs),
    .RESET_B(net1658),
    .D(net1751),
    .Q_N(\i_ibex/load_store_unit_i/_0451_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[16]_reg  (.RESET_B(net1658),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0051_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [16]),
    .Q_N(\i_ibex/load_store_unit_i/_0450_ ),
    .CLK(clknet_leaf_129_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[17]_reg  (.RESET_B(net1580),
    .VSS(VSS),
    .VDD(VDD),
    .D(net1726),
    .Q(\i_ibex/load_store_unit_i/rdata_q [17]),
    .Q_N(\i_ibex/load_store_unit_i/_0449_ ),
    .CLK(clknet_leaf_132_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[18]_reg  (.RESET_B(net1658),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0053_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [18]),
    .Q_N(\i_ibex/load_store_unit_i/_0448_ ),
    .CLK(clknet_leaf_129_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[19]_reg  (.RESET_B(net1581),
    .VSS(VSS),
    .VDD(VDD),
    .D(net1721),
    .Q(\i_ibex/load_store_unit_i/rdata_q [19]),
    .Q_N(\i_ibex/load_store_unit_i/_0447_ ),
    .CLK(clknet_leaf_130_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[1]_reg  (.CLK(clknet_leaf_132_clk_i_regs),
    .RESET_B(net1580),
    .D(net1747),
    .Q_N(\i_ibex/load_store_unit_i/_0446_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[20]_reg  (.RESET_B(net1659),
    .VSS(VSS),
    .VDD(VDD),
    .D(net1695),
    .Q(\i_ibex/load_store_unit_i/rdata_q [20]),
    .Q_N(\i_ibex/load_store_unit_i/_0445_ ),
    .CLK(clknet_leaf_134_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[21]_reg  (.RESET_B(net1659),
    .VSS(VSS),
    .VDD(VDD),
    .D(net1730),
    .Q(\i_ibex/load_store_unit_i/rdata_q [21]),
    .Q_N(\i_ibex/load_store_unit_i/_0444_ ),
    .CLK(clknet_leaf_130_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[22]_reg  (.RESET_B(net1580),
    .VSS(VSS),
    .VDD(VDD),
    .D(net1740),
    .Q(\i_ibex/load_store_unit_i/rdata_q [22]),
    .Q_N(\i_ibex/load_store_unit_i/_0443_ ),
    .CLK(clknet_leaf_133_clk_i_regs));
 sg13g2_dfrbp_2 \i_ibex/load_store_unit_i/rdata_q[23]_reg  (.RESET_B(net1658),
    .VSS(VSS),
    .VDD(VDD),
    .D(\i_ibex/load_store_unit_i/_0059_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [23]),
    .Q_N(\i_ibex/load_store_unit_i/_0442_ ),
    .CLK(clknet_leaf_135_clk_i_regs));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[2]_reg  (.CLK(clknet_leaf_130_clk_i_regs),
    .RESET_B(net1580),
    .D(net1737),
    .Q_N(\i_ibex/load_store_unit_i/_0441_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[3]_reg  (.CLK(clknet_leaf_132_clk_i_regs),
    .RESET_B(net1659),
    .D(net1734),
    .Q_N(\i_ibex/load_store_unit_i/_0440_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[4]_reg  (.CLK(clknet_leaf_130_clk_i_regs),
    .RESET_B(net1581),
    .D(net1743),
    .Q_N(\i_ibex/load_store_unit_i/_0439_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[5]_reg  (.CLK(clknet_leaf_130_clk_i_regs),
    .RESET_B(net1659),
    .D(net1714),
    .Q_N(\i_ibex/load_store_unit_i/_0438_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[6]_reg  (.CLK(clknet_leaf_133_clk_i_regs),
    .RESET_B(net1580),
    .D(net1716),
    .Q_N(\i_ibex/load_store_unit_i/_0437_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[7]_reg  (.CLK(clknet_leaf_128_clk_i_regs),
    .RESET_B(net1658),
    .D(net1753),
    .Q_N(\i_ibex/load_store_unit_i/_0436_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[8]_reg  (.CLK(clknet_leaf_128_clk_i_regs),
    .RESET_B(net1658),
    .D(net1749),
    .Q_N(\i_ibex/load_store_unit_i/_0435_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \i_ibex/load_store_unit_i/rdata_q[9]_reg  (.CLK(clknet_leaf_133_clk_i_regs),
    .RESET_B(net1580),
    .D(net1723),
    .Q_N(\i_ibex/load_store_unit_i/_0434_ ),
    .Q(\i_ibex/load_store_unit_i/rdata_q [9]),
    .VDD(VDD),
    .VSS(VSS));
 cve2_register_file_ff \i_ibex/register_file_i  (.VDD(VDD),
    .VSS(VSS),
    .clk_i(clknet_1_0__leaf_clk_i),
    .rst_ni(net1669),
    .test_en_i(test_enable_i),
    .we_a_i(\i_ibex/rf_we_wb ),
    .raddr_a_i({\i_ibex/id_stage_i/zimm_rs1_type [4],
    \i_ibex/id_stage_i/zimm_rs1_type [3],
    net765,
    net767,
    net769}),
    .raddr_b_i({net753,
    \i_ibex/id_stage_i/imm_u_type [23],
    net756,
    net760,
    net764}),
    .rdata_a_o({\i_ibex/rf_rdata_a [31],
    \i_ibex/rf_rdata_a [30],
    \i_ibex/rf_rdata_a [29],
    \i_ibex/rf_rdata_a [28],
    \i_ibex/rf_rdata_a [27],
    \i_ibex/rf_rdata_a [26],
    \i_ibex/rf_rdata_a [25],
    \i_ibex/rf_rdata_a [24],
    \i_ibex/rf_rdata_a [23],
    \i_ibex/rf_rdata_a [22],
    \i_ibex/rf_rdata_a [21],
    \i_ibex/rf_rdata_a [20],
    \i_ibex/rf_rdata_a [19],
    \i_ibex/rf_rdata_a [18],
    \i_ibex/rf_rdata_a [17],
    \i_ibex/rf_rdata_a [16],
    \i_ibex/rf_rdata_a [15],
    \i_ibex/rf_rdata_a [14],
    \i_ibex/rf_rdata_a [13],
    \i_ibex/rf_rdata_a [12],
    \i_ibex/rf_rdata_a [11],
    \i_ibex/rf_rdata_a [10],
    \i_ibex/rf_rdata_a [9],
    \i_ibex/rf_rdata_a [8],
    \i_ibex/rf_rdata_a [7],
    \i_ibex/rf_rdata_a [6],
    \i_ibex/rf_rdata_a [5],
    \i_ibex/rf_rdata_a [4],
    \i_ibex/rf_rdata_a [3],
    \i_ibex/rf_rdata_a [2],
    \i_ibex/rf_rdata_a [1],
    \i_ibex/rf_rdata_a [0]}),
    .rdata_b_o({\i_ibex/rf_rdata_b [31],
    \i_ibex/rf_rdata_b [30],
    \i_ibex/rf_rdata_b [29],
    \i_ibex/rf_rdata_b [28],
    \i_ibex/rf_rdata_b [27],
    \i_ibex/rf_rdata_b [26],
    \i_ibex/rf_rdata_b [25],
    \i_ibex/rf_rdata_b [24],
    \i_ibex/rf_rdata_b [23],
    \i_ibex/rf_rdata_b [22],
    \i_ibex/rf_rdata_b [21],
    \i_ibex/rf_rdata_b [20],
    \i_ibex/rf_rdata_b [19],
    \i_ibex/rf_rdata_b [18],
    \i_ibex/rf_rdata_b [17],
    \i_ibex/rf_rdata_b [16],
    \i_ibex/rf_rdata_b [15],
    \i_ibex/rf_rdata_b [14],
    \i_ibex/rf_rdata_b [13],
    \i_ibex/rf_rdata_b [12],
    \i_ibex/rf_rdata_b [11],
    \i_ibex/rf_rdata_b [10],
    \i_ibex/rf_rdata_b [9],
    \i_ibex/rf_rdata_b [8],
    \i_ibex/rf_rdata_b [7],
    \i_ibex/rf_rdata_b [6],
    \i_ibex/rf_rdata_b [5],
    \i_ibex/rf_rdata_b [4],
    \i_ibex/rf_rdata_b [3],
    \i_ibex/rf_rdata_b [2],
    \i_ibex/rf_rdata_b [1],
    \i_ibex/rf_rdata_b [0]}),
    .waddr_a_i({\i_ibex/id_stage_i/imm_s_type [4],
    \i_ibex/id_stage_i/imm_s_type [3],
    \i_ibex/id_stage_i/imm_s_type [2],
    \i_ibex/id_stage_i/imm_s_type [1],
    \i_ibex/id_stage_i/imm_s_type [0]}),
    .wdata_a_i({\i_ibex/rf_wdata_wb [31],
    \i_ibex/rf_wdata_wb [30],
    \i_ibex/rf_wdata_wb [29],
    \i_ibex/rf_wdata_wb [28],
    \i_ibex/rf_wdata_wb [27],
    \i_ibex/rf_wdata_wb [26],
    \i_ibex/rf_wdata_wb [25],
    \i_ibex/rf_wdata_wb [24],
    \i_ibex/rf_wdata_wb [23],
    \i_ibex/rf_wdata_wb [22],
    \i_ibex/rf_wdata_wb [21],
    \i_ibex/rf_wdata_wb [20],
    \i_ibex/rf_wdata_wb [19],
    \i_ibex/rf_wdata_wb [18],
    \i_ibex/rf_wdata_wb [17],
    \i_ibex/rf_wdata_wb [16],
    \i_ibex/rf_wdata_wb [15],
    \i_ibex/rf_wdata_wb [14],
    \i_ibex/rf_wdata_wb [13],
    \i_ibex/rf_wdata_wb [12],
    \i_ibex/rf_wdata_wb [11],
    \i_ibex/rf_wdata_wb [10],
    \i_ibex/rf_wdata_wb [9],
    \i_ibex/rf_wdata_wb [8],
    \i_ibex/rf_wdata_wb [7],
    \i_ibex/rf_wdata_wb [6],
    \i_ibex/rf_wdata_wb [5],
    \i_ibex/rf_wdata_wb [4],
    \i_ibex/rf_wdata_wb [3],
    \i_ibex/rf_wdata_wb [2],
    \i_ibex/rf_wdata_wb [1],
    \i_ibex/rf_wdata_wb [0]}));
 sg13g2_nand2_2 \i_ibex/wb_i/_040_  (.Y(\i_ibex/wb_i/_000_ ),
    .A(\i_ibex/lsu_resp_valid ),
    .B(\i_ibex/lsu_resp_err ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 \i_ibex/wb_i/_041_  (.X(\i_ibex/perf_instr_ret_wb ),
    .A(\i_ibex/instr_perf_count_id ),
    .B(\i_ibex/instr_id_done ),
    .C(\i_ibex/wb_i/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 \i_ibex/wb_i/_042_  (.A(\i_ibex/instr_perf_count_id ),
    .B(\i_ibex/instr_id_done ),
    .C(\i_ibex/instr_is_compressed_id ),
    .D(\i_ibex/wb_i/_000_ ),
    .X(\i_ibex/perf_instr_ret_compressed_wb ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout387 (.X(net387),
    .A(net389),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(net389),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_046_  (.Y(\i_ibex/wb_i/_004_ ),
    .B1(net1392),
    .B2(\i_ibex/rf_wdata_lsu [31]),
    .A2(\i_ibex/rf_wdata_id [31]),
    .A1(net969),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_047_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [31]),
    .A(\i_ibex/wb_i/_004_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_048_  (.Y(\i_ibex/wb_i/_005_ ),
    .B1(net1393),
    .B2(\i_ibex/rf_wdata_lsu [30]),
    .A2(\i_ibex/rf_wdata_id [30]),
    .A1(net970),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_049_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [30]),
    .A(\i_ibex/wb_i/_005_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_050_  (.Y(\i_ibex/wb_i/_006_ ),
    .B1(net1392),
    .B2(\i_ibex/rf_wdata_lsu [21]),
    .A2(\i_ibex/rf_wdata_id [21]),
    .A1(net969),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_051_  (.Y(\i_ibex/rf_wdata_wb [21]),
    .A(\i_ibex/wb_i/_006_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_052_  (.Y(\i_ibex/wb_i/_007_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [20]),
    .A2(\i_ibex/rf_wdata_id [20]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 \i_ibex/wb_i/_053_  (.A(\i_ibex/wb_i/_007_ ),
    .Y(\i_ibex/rf_wdata_wb [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_054_  (.Y(\i_ibex/wb_i/_008_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [19]),
    .A2(\i_ibex/rf_wdata_id [19]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_055_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [19]),
    .A(\i_ibex/wb_i/_008_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_056_  (.Y(\i_ibex/wb_i/_009_ ),
    .B1(net1392),
    .B2(\i_ibex/rf_wdata_lsu [18]),
    .A2(\i_ibex/rf_wdata_id [18]),
    .A1(net969),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_057_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [18]),
    .A(\i_ibex/wb_i/_009_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_058_  (.Y(\i_ibex/wb_i/_010_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [17]),
    .A2(\i_ibex/rf_wdata_id [17]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_059_  (.Y(\i_ibex/rf_wdata_wb [17]),
    .A(\i_ibex/wb_i/_010_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_060_  (.Y(\i_ibex/wb_i/_011_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [16]),
    .A2(\i_ibex/rf_wdata_id [16]),
    .A1(net969),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_061_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [16]),
    .A(\i_ibex/wb_i/_011_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_062_  (.Y(\i_ibex/wb_i/_012_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [15]),
    .A2(\i_ibex/rf_wdata_id [15]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_063_  (.Y(\i_ibex/rf_wdata_wb [15]),
    .A(\i_ibex/wb_i/_012_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(net389),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_065_  (.Y(\i_ibex/wb_i/_014_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [14]),
    .A2(\i_ibex/rf_wdata_id [14]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_066_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [14]),
    .A(\i_ibex/wb_i/_014_ ),
    .VSS(VSS));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(net389),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_068_  (.Y(\i_ibex/wb_i/_016_ ),
    .B1(net1390),
    .B2(\i_ibex/rf_wdata_lsu [13]),
    .A2(\i_ibex/rf_wdata_id [13]),
    .A1(net967),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_069_  (.Y(\i_ibex/rf_wdata_wb [13]),
    .A(\i_ibex/wb_i/_016_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_070_  (.Y(\i_ibex/wb_i/_017_ ),
    .B1(net1389),
    .B2(\i_ibex/rf_wdata_lsu [12]),
    .A2(\i_ibex/rf_wdata_id [12]),
    .A1(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_071_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [12]),
    .A(\i_ibex/wb_i/_017_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_072_  (.Y(\i_ibex/wb_i/_018_ ),
    .B1(net1390),
    .B2(\i_ibex/rf_wdata_lsu [29]),
    .A2(\i_ibex/rf_wdata_id [29]),
    .A1(net967),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_073_  (.Y(\i_ibex/rf_wdata_wb [29]),
    .A(\i_ibex/wb_i/_018_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_074_  (.Y(\i_ibex/wb_i/_019_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [11]),
    .A2(\i_ibex/rf_wdata_id [11]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_075_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [11]),
    .A(\i_ibex/wb_i/_019_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_076_  (.Y(\i_ibex/wb_i/_020_ ),
    .B1(net1389),
    .B2(\i_ibex/rf_wdata_lsu [10]),
    .A2(\i_ibex/rf_wdata_id [10]),
    .A1(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_077_  (.Y(\i_ibex/rf_wdata_wb [10]),
    .A(\i_ibex/wb_i/_020_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_078_  (.Y(\i_ibex/wb_i/_021_ ),
    .B1(net1390),
    .B2(\i_ibex/rf_wdata_lsu [9]),
    .A2(\i_ibex/rf_wdata_id [9]),
    .A1(net967),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_079_  (.Y(\i_ibex/rf_wdata_wb [9]),
    .A(\i_ibex/wb_i/_021_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_080_  (.Y(\i_ibex/wb_i/_022_ ),
    .B1(net1389),
    .B2(\i_ibex/rf_wdata_lsu [8]),
    .A2(\i_ibex/rf_wdata_id [8]),
    .A1(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_081_  (.Y(\i_ibex/rf_wdata_wb [8]),
    .A(\i_ibex/wb_i/_022_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_082_  (.Y(\i_ibex/wb_i/_023_ ),
    .B1(net1389),
    .B2(\i_ibex/rf_wdata_lsu [7]),
    .A2(\i_ibex/rf_wdata_id [7]),
    .A1(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_083_  (.Y(\i_ibex/rf_wdata_wb [7]),
    .A(\i_ibex/wb_i/_023_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_084_  (.Y(\i_ibex/wb_i/_024_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [6]),
    .A2(\i_ibex/rf_wdata_id [6]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_085_  (.Y(\i_ibex/rf_wdata_wb [6]),
    .A(\i_ibex/wb_i/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 fanout383 (.X(net383),
    .A(net389),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_087_  (.Y(\i_ibex/wb_i/_026_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [5]),
    .A2(\i_ibex/rf_wdata_id [5]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_088_  (.Y(\i_ibex/rf_wdata_wb [5]),
    .A(\i_ibex/wb_i/_026_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 max_cap382 (.X(net382),
    .A(net845),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_090_  (.Y(\i_ibex/wb_i/_028_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [4]),
    .A2(\i_ibex/rf_wdata_id [4]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_091_  (.Y(\i_ibex/rf_wdata_wb [4]),
    .A(\i_ibex/wb_i/_028_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_092_  (.Y(\i_ibex/wb_i/_029_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [3]),
    .A2(\i_ibex/rf_wdata_id [3]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_093_  (.Y(\i_ibex/rf_wdata_wb [3]),
    .A(\i_ibex/wb_i/_029_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_094_  (.Y(\i_ibex/wb_i/_030_ ),
    .B1(net1389),
    .B2(\i_ibex/rf_wdata_lsu [2]),
    .A2(\i_ibex/rf_wdata_id [2]),
    .A1(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_095_  (.Y(\i_ibex/rf_wdata_wb [2]),
    .A(\i_ibex/wb_i/_030_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_096_  (.Y(\i_ibex/wb_i/_031_ ),
    .B1(net1390),
    .B2(\i_ibex/rf_wdata_lsu [28]),
    .A2(\i_ibex/rf_wdata_id [28]),
    .A1(net967),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_097_  (.Y(\i_ibex/rf_wdata_wb [28]),
    .A(\i_ibex/wb_i/_031_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_098_  (.Y(\i_ibex/wb_i/_032_ ),
    .B1(net1388),
    .B2(\i_ibex/rf_wdata_lsu [1]),
    .A2(\i_ibex/rf_wdata_id [1]),
    .A1(net965),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_099_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [1]),
    .A(\i_ibex/wb_i/_032_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_100_  (.Y(\i_ibex/wb_i/_033_ ),
    .B1(net1389),
    .B2(\i_ibex/rf_wdata_lsu [0]),
    .A2(\i_ibex/rf_wdata_id [0]),
    .A1(net966),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_101_  (.Y(\i_ibex/rf_wdata_wb [0]),
    .A(\i_ibex/wb_i/_033_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_102_  (.Y(\i_ibex/wb_i/_034_ ),
    .B1(net1390),
    .B2(\i_ibex/rf_wdata_lsu [27]),
    .A2(\i_ibex/rf_wdata_id [27]),
    .A1(net967),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 \i_ibex/wb_i/_103_  (.A(\i_ibex/wb_i/_034_ ),
    .Y(\i_ibex/rf_wdata_wb [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_104_  (.Y(\i_ibex/wb_i/_035_ ),
    .B1(net1392),
    .B2(\i_ibex/rf_wdata_lsu [26]),
    .A2(\i_ibex/rf_wdata_id [26]),
    .A1(net969),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_105_  (.Y(\i_ibex/rf_wdata_wb [26]),
    .A(\i_ibex/wb_i/_035_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_106_  (.Y(\i_ibex/wb_i/_036_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [25]),
    .A2(\i_ibex/rf_wdata_id [25]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_107_  (.Y(\i_ibex/rf_wdata_wb [25]),
    .A(\i_ibex/wb_i/_036_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_108_  (.Y(\i_ibex/wb_i/_037_ ),
    .B1(net1392),
    .B2(\i_ibex/rf_wdata_lsu [24]),
    .A2(\i_ibex/rf_wdata_id [24]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 \i_ibex/wb_i/_109_  (.VDD(VDD),
    .Y(\i_ibex/rf_wdata_wb [24]),
    .A(\i_ibex/wb_i/_037_ ),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_110_  (.Y(\i_ibex/wb_i/_038_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [23]),
    .A2(\i_ibex/rf_wdata_id [23]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 \i_ibex/wb_i/_111_  (.Y(\i_ibex/rf_wdata_wb [23]),
    .A(\i_ibex/wb_i/_038_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 \i_ibex/wb_i/_112_  (.Y(\i_ibex/wb_i/_039_ ),
    .B1(net1391),
    .B2(\i_ibex/rf_wdata_lsu [22]),
    .A2(\i_ibex/rf_wdata_id [22]),
    .A1(net968),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 \i_ibex/wb_i/_113_  (.A(\i_ibex/wb_i/_039_ ),
    .Y(\i_ibex/rf_wdata_wb [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 \i_ibex/wb_i/_114_  (.VSS(VSS),
    .VDD(VDD),
    .X(\i_ibex/rf_we_wb ),
    .B(net1388),
    .A(net965));
 sg13g2_tielo \i_ibex/cs_registers_i/_1255__1  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net1));
 sg13g2_tielo \i_ibex/cs_registers_i/_1305__2  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net2));
 sg13g2_tielo \i_ibex/cs_registers_i/_1335__3  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net3));
 sg13g2_tielo \i_ibex/cs_registers_i/_1367__4  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net4));
 sg13g2_tielo \i_ibex/cs_registers_i/_1393__5  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net5));
 sg13g2_tielo \i_ibex/cs_registers_i/_1421__6  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net6));
 sg13g2_tielo \i_ibex/cs_registers_i/_1430__7  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net7));
 sg13g2_tielo \i_ibex/cs_registers_i/_1457__8  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net8));
 sg13g2_tielo \i_ibex/cs_registers_i/_1483__9  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net9));
 sg13g2_tielo \i_ibex/cs_registers_i/_1496__10  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net10));
 sg13g2_tielo \i_ibex/cs_registers_i/_1518__11  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net11));
 sg13g2_tielo \i_ibex/cs_registers_i/_1533__12  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net12));
 sg13g2_tielo \i_ibex/cs_registers_i/_1555__13  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net13));
 sg13g2_tielo \i_ibex/cs_registers_i/_1579__14  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net14));
 sg13g2_tielo \i_ibex/cs_registers_i/_1596__15  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net15));
 sg13g2_tielo \i_ibex/cs_registers_i/_1627__16  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net16));
 sg13g2_tielo \i_ibex/cs_registers_i/_1645__17  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net17));
 sg13g2_tielo \i_ibex/cs_registers_i/_1664__18  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net18));
 sg13g2_tielo \i_ibex/cs_registers_i/_1678__19  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net19));
 sg13g2_tielo \i_ibex/cs_registers_i/_1704__20  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net20));
 sg13g2_tielo \i_ibex/cs_registers_i/_1730__21  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net21));
 sg13g2_tielo \i_ibex/cs_registers_i/_1732__22  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net22));
 sg13g2_tielo \i_ibex/cs_registers_i/_1758__23  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net23));
 sg13g2_tielo \i_ibex/cs_registers_i/_1784__24  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net24));
 sg13g2_tielo \i_ibex/cs_registers_i/_1799__25  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net25));
 sg13g2_tielo \i_ibex/cs_registers_i/_1824__26  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net26));
 sg13g2_tielo \i_ibex/cs_registers_i/_1841__27  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net27));
 sg13g2_tielo \i_ibex/cs_registers_i/_1846__28  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net28));
 sg13g2_tielo \i_ibex/cs_registers_i/_1882__29  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net29));
 sg13g2_tielo \i_ibex/cs_registers_i/_1895__30  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net30));
 sg13g2_tielo \i_ibex/cs_registers_i/_1917__31  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net31));
 sg13g2_tielo \i_ibex/cs_registers_i/_1939__32  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net32));
 sg13g2_tielo \i_ibex/cs_registers_i/_1961__33  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net33));
 sg13g2_tielo \i_ibex/cs_registers_i/_1983__34  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net34));
 sg13g2_tielo \i_ibex/cs_registers_i/_2192__35  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net35));
 sg13g2_tielo \i_ibex/cs_registers_i/_2212__36  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net36));
 sg13g2_tielo \i_ibex/id_stage_i/controller_i/_662__37  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net37));
 sg13g2_tielo \i_ibex/id_stage_i/controller_i/_671__38  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net38));
 sg13g2_tielo \i_ibex/id_stage_i/controller_i/_783__39  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net39));
 sg13g2_tielo \i_ibex/id_stage_i/controller_i/_794__40  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net40));
 sg13g2_tielo \i_ibex/id_stage_i/controller_i/_858__41  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net41));
 sg13g2_tielo \i_ibex/if_stage_i/_736__43  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net43));
 sg13g2_tielo \i_ibex/if_stage_i/_740__44  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net44));
 sg13g2_tielo \i_ibex/load_store_unit_i/_0969__45  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net45));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_085__47  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net47));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_097__48  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net48));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_100__49  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net49));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_101__50  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net50));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_102__51  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net51));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_103__52  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net52));
 sg13g2_tielo \i_ibex/cs_registers_i/u_mtvec_csr/_104__53  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net53));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1475__73  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net73));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1477__74  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net74));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1477__75  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net75));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1480__76  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net76));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1484__77  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net77));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1492__78  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net78));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1493__79  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net79));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1497__80  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net80));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1499__81  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net81));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1499__82  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net82));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1505__83  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net83));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1506__84  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net84));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1519__85  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net85));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1523__86  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net86));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1523__87  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net87));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1527__88  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net88));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1527__89  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net89));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1532__90  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net90));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1536__91  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net91));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1540__92  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net92));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1540__93  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net93));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1545__94  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net94));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1545__95  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net95));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1546__96  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net96));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1546__97  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net97));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1550__98  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net98));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1550__99  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net99));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1555__100  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net100));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1557__101  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net101));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1558__102  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net102));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1564__103  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net103));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1565__104  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net104));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1565__105  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net105));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1566__106  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net106));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1566__107  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net107));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1570__108  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net108));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1570__109  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net109));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1577__110  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net110));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1577__111  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net111));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1585__112  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net112));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1586__113  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net113));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1595__114  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net114));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1595__115  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net115));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1596__116  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net116));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1596__117  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net117));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1602__118  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net118));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1603__119  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net119));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1610__120  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net120));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1611__121  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net121));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1621__122  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net122));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1622__123  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net123));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1626__124  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net124));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1627__125  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net125));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1634__126  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net126));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1635__127  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net127));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1642__128  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net128));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1643__129  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net129));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1650__130  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net130));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1652__131  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net131));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1661__132  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net132));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1664__133  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net133));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1665__134  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net134));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1668__135  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net135));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1668__136  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net136));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1670__137  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net137));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1670__138  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net138));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1672__139  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net139));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1679__140  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net140));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1680__141  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net141));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1683__142  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net142));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1696__143  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net143));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1696__144  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net144));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1700__145  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net145));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1703__146  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net146));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1705__147  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net147));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1705__148  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net148));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1710__149  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net149));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1712__150  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net150));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1712__151  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net151));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1714__152  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net152));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1716__153  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net153));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1716__154  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net154));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1719__155  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net155));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1719__156  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net156));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1725__157  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net157));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1725__158  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net158));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1730__159  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net159));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1731__160  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net160));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1741__161  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net161));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1741__162  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net162));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1742__163  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net163));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1742__164  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net164));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1747__165  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net165));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1748__166  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net166));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1756__167  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net167));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1759__168  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net168));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1764__169  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net169));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1766__170  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net170));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1766__171  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net171));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1770__172  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net172));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1772__173  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net173));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1772__174  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net174));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1777__175  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net175));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1778__176  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net176));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1778__177  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net177));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1784__178  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net178));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1784__179  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net179));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1787__180  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net180));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1790__181  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net181));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1790__182  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net182));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1793__183  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net183));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1802__184  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net184));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1802__185  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net185));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1804__186  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net186));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1804__187  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net187));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1807__188  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net188));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1810__189  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net189));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1811__190  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net190));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1811__191  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net191));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1820__192  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net192));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1820__193  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net193));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1823__194  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net194));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1825__195  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net195));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1825__196  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net196));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1829__197  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net197));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1829__198  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net198));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1834__199  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net199));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1834__200  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net200));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1836__201  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net201));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1838__202  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net202));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1838__203  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net203));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1840__204  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net204));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1842__205  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net205));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1842__206  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net206));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1846__207  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net207));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1847__208  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net208));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1847__209  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net209));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1857__210  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net210));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1858__211  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net211));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1865__212  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net212));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1866__213  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net213));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1875__214  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net214));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1876__215  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net215));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1883__216  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net216));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1884__217  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net217));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1889__218  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net218));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1891__219  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net219));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1892__220  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net220));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1893__221  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net221));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1893__222  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net222));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1901__223  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net223));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1903__224  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net224));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1903__225  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net225));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1907__226  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net226));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1907__227  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net227));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1912__228  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net228));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1912__229  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net229));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1916__230  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net230));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1918__231  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net231));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1918__232  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net232));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1924__233  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net233));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1926__234  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net234));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1931__235  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net235));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1933__236  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net236));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1950__237  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net237));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1950__238  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net238));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2018__239  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net239));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2020__240  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net240));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2029__241  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net241));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2031__242  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net242));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2036__243  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net243));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2037__244  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net244));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2038__245  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net245));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2038__246  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net246));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2039__247  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net247));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2042__248  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net248));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2045__249  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net249));
 sg13g2_tielo \i_ibex/id_stage_i/_1199__250  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net250));
 sg13g2_tielo \i_ibex/id_stage_i/_1200__251  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net251));
 sg13g2_tielo \i_ibex/id_stage_i/_1240__252  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net252));
 sg13g2_tielo \i_ibex/id_stage_i/_1241__253  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net253));
 sg13g2_tielo \i_ibex/ex_block_i/_1__255  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net255));
 sg13g2_tielo \i_ibex/id_stage_i/_1170__256  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net256));
 sg13g2_tielo \i_ibex/id_stage_i/_1172__257  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net257));
 sg13g2_tielo \i_ibex/id_stage_i/_1173__258  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net258));
 sg13g2_tielo \i_ibex/id_stage_i/_1174__259  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net259));
 sg13g2_tielo \i_ibex/id_stage_i/_1175__260  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net260));
 sg13g2_tielo \i_ibex/id_stage_i/_1176__261  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net261));
 sg13g2_tielo \i_ibex/id_stage_i/_1177__262  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net262));
 sg13g2_tielo \i_ibex/id_stage_i/_1178__263  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net263));
 sg13g2_tielo \i_ibex/id_stage_i/_1179__264  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net264));
 sg13g2_tielo \i_ibex/id_stage_i/_1180__265  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net265));
 sg13g2_tielo \i_ibex/id_stage_i/_1181__266  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net266));
 sg13g2_tielo \i_ibex/id_stage_i/_1183__267  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net267));
 sg13g2_tielo \i_ibex/id_stage_i/_1184__268  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net268));
 sg13g2_tielo \i_ibex/id_stage_i/_1185__269  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net269));
 sg13g2_tielo \i_ibex/id_stage_i/_1186__270  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net270));
 sg13g2_tielo \i_ibex/id_stage_i/_1187__271  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net271));
 sg13g2_tielo \i_ibex/id_stage_i/_1188__272  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net272));
 sg13g2_tielo \i_ibex/id_stage_i/_1189__273  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net273));
 sg13g2_tielo \i_ibex/id_stage_i/_1190__274  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net274));
 sg13g2_tielo \i_ibex/id_stage_i/_1191__275  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net275));
 sg13g2_tielo \i_ibex/id_stage_i/_1192__276  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net276));
 sg13g2_tielo \i_ibex/id_stage_i/_1194__277  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net277));
 sg13g2_tielo \i_ibex/id_stage_i/_1195__278  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net278));
 sg13g2_tielo \i_ibex/id_stage_i/_1196__279  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net279));
 sg13g2_tielo \i_ibex/id_stage_i/_1197__280  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net280));
 sg13g2_tielo \i_ibex/id_stage_i/_1198__281  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net281));
 sg13g2_tielo \i_ibex/id_stage_i/_1201__282  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net282));
 sg13g2_tielo \i_ibex/id_stage_i/_1203__283  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net283));
 sg13g2_tielo \i_ibex/id_stage_i/_1204__284  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net284));
 sg13g2_tielo \i_ibex/id_stage_i/_1205__285  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net285));
 sg13g2_tielo \i_ibex/id_stage_i/_1206__286  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net286));
 sg13g2_tielo \i_ibex/id_stage_i/_1207__287  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net287));
 sg13g2_tielo \i_ibex/id_stage_i/_1208__288  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net288));
 sg13g2_tielo \i_ibex/id_stage_i/_1209__289  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net289));
 sg13g2_tielo \i_ibex/id_stage_i/_1210__290  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net290));
 sg13g2_tielo \i_ibex/id_stage_i/_1211__291  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net291));
 sg13g2_tielo \i_ibex/id_stage_i/_1212__292  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net292));
 sg13g2_tielo \i_ibex/id_stage_i/_1213__293  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net293));
 sg13g2_tielo \i_ibex/id_stage_i/_1215__294  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net294));
 sg13g2_tielo \i_ibex/id_stage_i/_1216__295  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net295));
 sg13g2_tielo \i_ibex/id_stage_i/_1217__296  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net296));
 sg13g2_tielo \i_ibex/id_stage_i/_1218__297  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net297));
 sg13g2_tielo \i_ibex/id_stage_i/_1219__298  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net298));
 sg13g2_tielo \i_ibex/id_stage_i/_1220__299  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net299));
 sg13g2_tielo \i_ibex/id_stage_i/_1221__300  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net300));
 sg13g2_tielo \i_ibex/id_stage_i/_1222__301  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net301));
 sg13g2_tielo \i_ibex/id_stage_i/_1223__302  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net302));
 sg13g2_tielo \i_ibex/id_stage_i/_1224__303  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net303));
 sg13g2_tielo \i_ibex/id_stage_i/_1225__304  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net304));
 sg13g2_tielo \i_ibex/id_stage_i/_1227__305  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net305));
 sg13g2_tielo \i_ibex/id_stage_i/_1228__306  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net306));
 sg13g2_tielo \i_ibex/id_stage_i/_1229__307  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net307));
 sg13g2_tielo \i_ibex/id_stage_i/_1230__308  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net308));
 sg13g2_tielo \i_ibex/id_stage_i/_1231__309  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net309));
 sg13g2_tielo \i_ibex/id_stage_i/_1232__310  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net310));
 sg13g2_tielo \i_ibex/id_stage_i/_1233__311  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net311));
 sg13g2_tielo \i_ibex/id_stage_i/_1234__312  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net312));
 sg13g2_tielo \i_ibex/id_stage_i/_1235__313  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net313));
 sg13g2_tielo \i_ibex/id_stage_i/_1236__314  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net314));
 sg13g2_tielo \i_ibex/id_stage_i/_1237__315  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net315));
 sg13g2_tielo \i_ibex/id_stage_i/_1238__316  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net316));
 sg13g2_tielo \i_ibex/id_stage_i/_1239__317  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net317));
 sg13g2_tielo \i_ibex/id_stage_i/_1242__318  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net318));
 sg13g2_tielo \i_ibex/id_stage_i/_1243__319  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net319));
 sg13g2_tielo \i_ibex/id_stage_i/_1244__320  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net320));
 sg13g2_tielo \i_ibex/id_stage_i/_1245__321  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net321));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1369__323  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net323));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_1377__324  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net324));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2061__325  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net325));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2066__326  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net326));
 sg13g2_tielo \i_ibex/ex_block_i/alu_i/_2207__327  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net327));
 sg13g2_tielo \i_ibex/id_stage_i/_0645__328  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net328));
 sg13g2_tielo \i_ibex/id_stage_i/_0650__329  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net329));
 sg13g2_tielo \i_ibex/id_stage_i/_0655__330  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net330));
 sg13g2_tielo \i_ibex/id_stage_i/_0660__331  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net331));
 sg13g2_tielo \i_ibex/id_stage_i/_0665__332  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net332));
 sg13g2_tielo \i_ibex/id_stage_i/_0670__333  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net333));
 sg13g2_tielo \i_ibex/id_stage_i/_0676__334  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net334));
 sg13g2_tielo \i_ibex/id_stage_i/_0681__335  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net335));
 sg13g2_tielo \i_ibex/id_stage_i/_0686__336  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net336));
 sg13g2_tielo \i_ibex/id_stage_i/_0692__337  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net337));
 sg13g2_tielo \i_ibex/id_stage_i/_0702__338  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net338));
 sg13g2_tielo \i_ibex/id_stage_i/_0707__339  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net339));
 sg13g2_tielo \i_ibex/id_stage_i/_0712__340  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net340));
 sg13g2_tielo \i_ibex/id_stage_i/_0717__341  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net341));
 sg13g2_tielo \i_ibex/id_stage_i/_0722__342  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net342));
 sg13g2_tielo \i_ibex/id_stage_i/_0727__343  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net343));
 sg13g2_tielo \i_ibex/id_stage_i/_0733__344  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net344));
 sg13g2_tielo \i_ibex/id_stage_i/_0738__345  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net345));
 sg13g2_tielo \i_ibex/id_stage_i/_0743__346  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net346));
 sg13g2_tielo \i_ibex/id_stage_i/_0749__347  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net347));
 sg13g2_tielo \i_ibex/id_stage_i/_0774__348  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net348));
 sg13g2_tielo \i_ibex/id_stage_i/_0789__349  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net349));
 sg13g2_tielo \i_ibex/id_stage_i/_0794__350  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net350));
 sg13g2_tielo \i_ibex/id_stage_i/_0799__351  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net351));
 sg13g2_tielo \i_ibex/id_stage_i/_0804__352  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net352));
 sg13g2_tielo \i_ibex/id_stage_i/_0809__353  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net353));
 sg13g2_tielo \i_ibex/id_stage_i/_0814__354  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net354));
 sg13g2_tielo \i_ibex/id_stage_i/_0954__355  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net355));
 sg13g2_tielo \i_ibex/id_stage_i/_0962__356  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net356));
 sg13g2_tielo \i_ibex/id_stage_i/_0970__357  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net357));
 sg13g2_tielo \i_ibex/id_stage_i/_0979__358  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net358));
 sg13g2_tielo \i_ibex/id_stage_i/_0988__359  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net359));
 sg13g2_tielo \i_ibex/id_stage_i/_0997__360  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net360));
 sg13g2_tielo \i_ibex/id_stage_i/_1006__361  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net361));
 sg13g2_tielo \i_ibex/id_stage_i/_1016__362  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net362));
 sg13g2_tielo \i_ibex/id_stage_i/_1026__363  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net363));
 sg13g2_tielo \i_ibex/id_stage_i/_1034__364  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net364));
 sg13g2_tielo \i_ibex/id_stage_i/_1058__365  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net365));
 sg13g2_tielo \i_ibex/id_stage_i/_1065__366  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net366));
 sg13g2_tielo \i_ibex/id_stage_i/_1066__367  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net367));
 sg13g2_tielo \i_ibex/id_stage_i/_1069__368  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net368));
 sg13g2_tielo \i_ibex/id_stage_i/_1135__369  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net369));
 sg13g2_tielo \i_ibex/id_stage_i/_1135__370  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net370));
 sg13g2_tielo \i_ibex/id_stage_i/_1137__371  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net371));
 sg13g2_tielo \i_ibex/id_stage_i/_1160__372  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net372));
 sg13g2_tielo \i_ibex/id_stage_i/_1162__373  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net373));
 sg13g2_tielo \i_ibex/id_stage_i/_1162__374  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net374));
 sg13g2_tielo \i_ibex/id_stage_i/_1164__375  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net375));
 sg13g2_tielo \i_ibex/id_stage_i/_1254__376  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net376));
 sg13g2_tielo \i_ibex/id_stage_i/_1299__377  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net377));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(net1052),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout1052 (.A(\i_ibex/ex_block_i/alu_i/_0802_ ),
    .X(net1052),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1056),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1054 (.A(net1056),
    .X(net1054),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1055 (.A(net1056),
    .X(net1055),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(\i_ibex/cs_registers_i/_0952_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1058 (.X(net1058),
    .A(net1059),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(net1060),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1060 (.A(\i_ibex/cs_registers_i/_0952_ ),
    .X(net1060),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(\i_ibex/cs_registers_i/_0013_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(net1064),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1064),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1064 (.A(net1073),
    .X(net1064),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1065 (.A(net1066),
    .X(net1065),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1066 (.A(net1067),
    .X(net1066),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1067 (.A(net1073),
    .X(net1067),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1068 (.A(net1073),
    .X(net1068),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1069 (.A(net1070),
    .X(net1069),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1070 (.A(net1071),
    .X(net1070),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1071 (.A(net1072),
    .X(net1071),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1072 (.A(net1073),
    .X(net1072),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1073 (.A(net485),
    .X(net1073),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1076),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1076 (.A(net1078),
    .X(net1076),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1077 (.X(net1077),
    .A(net1078),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1079 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_181_ ),
    .X(net1079),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1084),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(net1082),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1082 (.A(net1083),
    .X(net1082),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1083 (.A(net1084),
    .X(net1083),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1084 (.A(\i_ibex/csr_mtvec_init ),
    .X(net1084),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1085 (.A(net1086),
    .X(net1085),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1086 (.A(net1087),
    .X(net1086),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1087 (.A(\i_ibex/ex_block_i/alu_i/_0103_ ),
    .X(net1087),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1088 (.A(net1089),
    .X(net1088),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(\i_ibex/csr_addr [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1090 (.A(net1092),
    .X(net1090),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1091 (.A(net1092),
    .X(net1091),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1092 (.A(\i_ibex/csr_addr [4]),
    .X(net1092),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1093 (.A(net1096),
    .X(net1093),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1094 (.A(net1095),
    .X(net1094),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1096 (.A(\i_ibex/csr_addr [6]),
    .X(net1096),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1097 (.A(net1098),
    .X(net1097),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1098 (.A(\i_ibex/csr_addr [7]),
    .X(net1098),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1099 (.X(net1099),
    .A(net1105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1100 (.A(net1105),
    .X(net1100),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1101 (.A(net1102),
    .X(net1101),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1102 (.A(net1103),
    .X(net1102),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1104 (.A(net1105),
    .X(net1104),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1105 (.A(\i_ibex/csr_addr [0]),
    .X(net1105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1106 (.A(\i_ibex/csr_addr [10]),
    .X(net1106),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1107 (.A(\i_ibex/alu_operand_b_ex [12]),
    .X(net1107),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1108 (.A(net1109),
    .X(net1108),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1109 (.A(net1110),
    .X(net1109),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1110 (.A(\i_ibex/ex_block_i/alu_i/_0072_ ),
    .X(net1110),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1111 (.A(net1112),
    .X(net1111),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1112 (.A(\i_ibex/ex_block_i/alu_i/_0072_ ),
    .X(net1112),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1113 (.A(\i_ibex/cs_registers_i/_0881_ ),
    .X(net1113),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1114 (.A(net1117),
    .X(net1114),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1115 (.A(net1117),
    .X(net1115),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1117 (.A(net1121),
    .X(net1117),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1118 (.A(net1120),
    .X(net1118),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1119 (.A(net1120),
    .X(net1119),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1120 (.A(net1121),
    .X(net1120),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1121 (.A(net523),
    .X(net1121),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1122 (.A(net1126),
    .X(net1122),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1123 (.A(net1126),
    .X(net1123),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1124 (.A(net1125),
    .X(net1124),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1125 (.A(net1126),
    .X(net1125),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(net524),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1127 (.A(net1128),
    .X(net1127),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1128 (.A(net1129),
    .X(net1128),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1129 (.A(net1132),
    .X(net1129),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1130 (.A(net1132),
    .X(net1130),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1131 (.A(net1132),
    .X(net1131),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1132 (.A(net525),
    .X(net1132),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1133 (.X(net1133),
    .A(net1137),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(net1137),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1135 (.X(net1135),
    .A(net1136),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1136 (.X(net1136),
    .A(net1137),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1137 (.A(\i_ibex/load_store_unit_i/_0098_ ),
    .X(net1137),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1138 (.X(net1138),
    .A(net1139),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1139 (.A(\i_ibex/pc_set ),
    .X(net1139),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(\i_ibex/pc_set ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1141 (.A(net1143),
    .X(net1141),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1142 (.A(net1143),
    .X(net1142),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1143 (.A(\i_ibex/ex_block_i/alu_i/_0152_ ),
    .X(net1143),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1144 (.A(net1145),
    .X(net1144),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1145 (.A(\i_ibex/ex_block_i/alu_i/_0152_ ),
    .X(net1145),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1146 (.A(net1147),
    .X(net1146),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1147 (.A(net1150),
    .X(net1147),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1148 (.A(net1149),
    .X(net1148),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(net1150),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1150 (.A(\i_ibex/ex_block_i/alu_i/_0066_ ),
    .X(net1150),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1151 (.A(\i_ibex/ex_block_i/alu_i/_1287_ ),
    .X(net1151),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1152 (.A(net1153),
    .X(net1152),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(\i_ibex/ex_block_i/alu_i/_0721_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1154 (.A(net1155),
    .X(net1154),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1155 (.A(\i_ibex/ex_block_i/alu_i/_0721_ ),
    .X(net1155),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(net1158),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1157 (.A(net1158),
    .X(net1157),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1158 (.A(net1159),
    .X(net1158),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(\i_ibex/ex_block_i/alu_i/_0670_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1160 (.A(net1163),
    .X(net1160),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1161 (.A(net1163),
    .X(net1161),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1162 (.A(net1163),
    .X(net1162),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1163 (.A(net1170),
    .X(net1163),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1164 (.A(net1170),
    .X(net1164),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1165 (.A(net1170),
    .X(net1165),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1166 (.A(net1168),
    .X(net1166),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1167 (.A(net1168),
    .X(net1167),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1168 (.A(net1169),
    .X(net1168),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1169 (.A(net1170),
    .X(net1169),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1170 (.A(\i_ibex/ex_block_i/alu_i/_0150_ ),
    .X(net1170),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1171 (.A(net1173),
    .X(net1171),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1172 (.A(net1173),
    .X(net1172),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1173 (.A(net1176),
    .X(net1173),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1174 (.A(net1175),
    .X(net1174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1175 (.A(net1176),
    .X(net1175),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1176 (.A(\i_ibex/ex_block_i/alu_i/_0149_ ),
    .X(net1176),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1177 (.A(net1178),
    .X(net1177),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1178 (.A(net1181),
    .X(net1178),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1179 (.A(net1180),
    .X(net1179),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(net1181),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1181 (.A(\i_ibex/ex_block_i/alu_i/_0069_ ),
    .X(net1181),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1182 (.X(net1182),
    .A(net1183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1183 (.A(net1184),
    .X(net1183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1184 (.A(net1187),
    .X(net1184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1185 (.A(net1186),
    .X(net1185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1186 (.A(net1187),
    .X(net1186),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1187 (.A(\i_ibex/if_stage_i/_093_ ),
    .X(net1187),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1188 (.A(net1192),
    .X(net1188),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1189 (.A(net1192),
    .X(net1189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1190 (.A(net1192),
    .X(net1190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1191 (.A(net1192),
    .X(net1191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1192 (.A(\i_ibex/id_stage_i/_0523_ ),
    .X(net1192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1193 (.A(net1195),
    .X(net1193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1194 (.A(net1195),
    .X(net1194),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1195 (.A(\i_ibex/id_stage_i/_0368_ ),
    .X(net1195),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1196 (.A(net1197),
    .X(net1196),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1197 (.A(\i_ibex/id_stage_i/_0368_ ),
    .X(net1197),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1198 (.X(net1198),
    .A(net1202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1199 (.A(net1202),
    .X(net1199),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1200 (.A(net1202),
    .X(net1200),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1201 (.A(net1202),
    .X(net1201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1202 (.A(net1205),
    .X(net1202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1203 (.X(net1203),
    .A(net1204),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1204 (.A(net1205),
    .X(net1204),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1205 (.A(\i_ibex/ex_block_i/alu_i/_0089_ ),
    .X(net1205),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1206 (.X(net1206),
    .A(net1208),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1207 (.A(net1208),
    .X(net1207),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1208 (.X(net1208),
    .A(net1211),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1209 (.X(net1209),
    .A(net1210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1210 (.X(net1210),
    .A(net1211),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1211 (.A(\i_ibex/ex_block_i/alu_i/_0076_ ),
    .X(net1211),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1212 (.A(net1213),
    .X(net1212),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net1217),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1214 (.A(net1217),
    .X(net1214),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1215 (.A(net1217),
    .X(net1215),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1216 (.A(net1217),
    .X(net1216),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1217 (.A(\i_ibex/ex_block_i/alu_i/_0070_ ),
    .X(net1217),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1218 (.A(net1221),
    .X(net1218),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1220 (.A(net1221),
    .X(net1220),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1221 (.X(net1221),
    .A(\i_ibex/if_stage_i/_112_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(net1223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1223 (.A(net1226),
    .X(net1223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1224 (.X(net1224),
    .A(net1225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1225 (.A(net1226),
    .X(net1225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1226 (.A(\i_ibex/if_stage_i/_111_ ),
    .X(net1226),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1227 (.A(\i_ibex/if_stage_i/_100_ ),
    .X(net1227),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1228 (.A(net1229),
    .X(net1228),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1229 (.A(net1230),
    .X(net1229),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1230 (.A(\i_ibex/if_stage_i/_100_ ),
    .X(net1230),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1231 (.A(\i_ibex/if_stage_i/_098_ ),
    .X(net1231),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1232 (.A(net1233),
    .X(net1232),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1233 (.A(net1234),
    .X(net1233),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1234 (.A(\i_ibex/if_stage_i/_098_ ),
    .X(net1234),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1235 (.A(net1236),
    .X(net1235),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1236 (.A(net1239),
    .X(net1236),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1237 (.A(net1238),
    .X(net1237),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1238 (.A(net1239),
    .X(net1238),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1239 (.A(\i_ibex/if_stage_i/_096_ ),
    .X(net1239),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1240 (.A(net1241),
    .X(net1240),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1241 (.A(\i_ibex/id_stage_i/_0537_ ),
    .X(net1241),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1242 (.A(net1243),
    .X(net1242),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1243 (.A(\i_ibex/id_stage_i/_0537_ ),
    .X(net1243),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1244 (.A(net1248),
    .X(net1244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1245 (.A(net1248),
    .X(net1245),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1246 (.A(net1248),
    .X(net1246),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1247 (.A(net1248),
    .X(net1247),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1248 (.A(\i_ibex/id_stage_i/_0530_ ),
    .X(net1248),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1249 (.A(net1253),
    .X(net1249),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1250 (.A(net1253),
    .X(net1250),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1251 (.A(net1253),
    .X(net1251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1252 (.A(net1253),
    .X(net1252),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1253 (.A(\i_ibex/id_stage_i/_0520_ ),
    .X(net1253),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1254 (.A(net1256),
    .X(net1254),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1255 (.A(net1256),
    .X(net1255),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1256 (.A(\i_ibex/id_stage_i/_0366_ ),
    .X(net1256),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1258 (.A(\i_ibex/id_stage_i/_0366_ ),
    .X(net1258),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1259 (.A(net1264),
    .X(net1259),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1260 (.A(net1264),
    .X(net1260),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1261 (.A(net1263),
    .X(net1261),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1262 (.A(net1264),
    .X(net1262),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1263 (.A(net1264),
    .X(net1263),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1264 (.A(\i_ibex/id_stage_i/_0361_ ),
    .X(net1264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1265 (.A(net1267),
    .X(net1265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1266 (.A(net1267),
    .X(net1266),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1267 (.A(net1268),
    .X(net1267),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1268 (.X(net1268),
    .A(\i_ibex/cs_registers_i/_0950_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1269 (.X(net1269),
    .A(net1270),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(net1271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1271 (.A(\i_ibex/cs_registers_i/_0950_ ),
    .X(net1271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1272 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_113_ ),
    .X(net1272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1273 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_045_ ),
    .X(net1273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1274 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_424_ ),
    .X(net1274),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1275 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_424_ ),
    .X(net1275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1276 (.A(net1277),
    .X(net1276),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1277 (.A(\i_ibex/load_store_unit_i/_0244_ ),
    .X(net1277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1278 (.A(net1279),
    .X(net1278),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1279 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_198_ ),
    .X(net1279),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1280 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_032_ ),
    .X(net1280),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1281 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_028_ ),
    .X(net1281),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1282 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_028_ ),
    .X(net1282),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1283 (.X(net1283),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_000_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1284 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_000_ ),
    .X(net1284),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1285 (.A(net1286),
    .X(net1285),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1286 (.A(net1287),
    .X(net1286),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1287 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_433_ ),
    .X(net1287),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1288 (.A(net1289),
    .X(net1288),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1289 (.A(\i_ibex/alu_operator_ex [0]),
    .X(net1289),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1290 (.A(\i_ibex/alu_operator_ex [2]),
    .X(net1290),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1291 (.A(\i_ibex/alu_operator_ex [2]),
    .X(net1291),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1292 (.A(net1293),
    .X(net1292),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1293 (.A(\i_ibex/alu_operator_ex [3]),
    .X(net1293),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1294 (.A(net1296),
    .X(net1294),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1295 (.A(net1296),
    .X(net1295),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1296 (.A(net1299),
    .X(net1296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1297 (.A(net1298),
    .X(net1297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1299 (.X(net1299),
    .A(\i_ibex/id_stage_i/alu_op_a_mux_sel_dec [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1300 (.A(net1301),
    .X(net1300),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1301 (.A(net1304),
    .X(net1301),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1302 (.A(net1303),
    .X(net1302),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1303 (.A(net1304),
    .X(net1303),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1304 (.A(\i_ibex/id_stage_i/alu_op_a_mux_sel_dec [1]),
    .X(net1304),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1305 (.X(net1305),
    .A(net1306),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1306 (.A(net1309),
    .X(net1306),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1307 (.A(net1308),
    .X(net1307),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1308 (.A(net1309),
    .X(net1308),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1309 (.A(net1315),
    .X(net1309),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1310 (.A(net1311),
    .X(net1310),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1311 (.A(net1313),
    .X(net1311),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1312 (.A(net1313),
    .X(net1312),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1313 (.A(net1315),
    .X(net1313),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1314 (.A(net1315),
    .X(net1314),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1315 (.A(\i_ibex/pc_mux_id [1]),
    .X(net1315),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1316 (.X(net1316),
    .A(net1320),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1317 (.A(net1320),
    .X(net1317),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1318 (.X(net1318),
    .A(net1320),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1319 (.A(net1320),
    .X(net1319),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1320 (.A(\i_ibex/load_store_unit_i/_0430_ ),
    .X(net1320),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1321 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/_083_ ),
    .X(net1321),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1322 (.X(net1322),
    .A(\i_ibex/if_stage_i/compressed_decoder_i/_024_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1323 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_019_ ),
    .X(net1323),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1324 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_019_ ),
    .X(net1324),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1325 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_414_ ),
    .X(net1325),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1326 (.A(\i_ibex/if_stage_i/compressed_decoder_i/_414_ ),
    .X(net1326),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1327 (.A(net1328),
    .X(net1327),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1328 (.A(net1331),
    .X(net1328),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1329 (.A(net1331),
    .X(net1329),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1330 (.A(net1331),
    .X(net1330),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1331 (.A(net1337),
    .X(net1331),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1332 (.A(net1333),
    .X(net1332),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1333 (.A(net1337),
    .X(net1333),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1334 (.A(net1336),
    .X(net1334),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1335 (.A(net1336),
    .X(net1335),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1336 (.A(net1337),
    .X(net1336),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1337 (.A(\i_ibex/id_stage_i/imm_b_mux_sel_dec [2]),
    .X(net1337),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1338 (.A(net1339),
    .X(net1338),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1339 (.A(net1342),
    .X(net1339),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1340 (.A(net1341),
    .X(net1340),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1341 (.A(net1342),
    .X(net1341),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1342 (.A(\i_ibex/exc_pc_mux_id [1]),
    .X(net1342),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1343 (.A(net1344),
    .X(net1343),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1344 (.A(net1346),
    .X(net1344),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1345 (.A(net1346),
    .X(net1345),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1346 (.A(net1349),
    .X(net1346),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1347 (.A(net1348),
    .X(net1347),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1348 (.A(net1349),
    .X(net1348),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1349 (.A(\i_ibex/if_stage_i/fetch_rdata [1]),
    .X(net1349),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1350 (.A(\i_ibex/if_stage_i/fetch_rdata [2]),
    .X(net1350),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1351 (.A(\i_ibex/if_stage_i/fetch_rdata [3]),
    .X(net1351),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1352 (.A(\i_ibex/if_stage_i/fetch_rdata [3]),
    .X(net1352),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1353 (.X(net1353),
    .A(\i_ibex/if_stage_i/fetch_rdata [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1354 (.A(\i_ibex/if_stage_i/fetch_rdata [7]),
    .X(net1354),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1355 (.A(\i_ibex/if_stage_i/fetch_rdata [7]),
    .X(net1355),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1356 (.A(net1357),
    .X(net1356),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1357 (.A(\i_ibex/if_stage_i/fetch_rdata [9]),
    .X(net1357),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1358 (.A(net1359),
    .X(net1358),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1359 (.A(\i_ibex/if_stage_i/fetch_rdata [10]),
    .X(net1359),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1360 (.X(net1360),
    .A(net1361),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1361 (.A(net1362),
    .X(net1361),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1362 (.X(net1362),
    .A(net1365),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1363 (.X(net1363),
    .A(net1364),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1364 (.A(net1365),
    .X(net1364),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1365 (.A(\i_ibex/id_stage_i/rf_wdata_sel ),
    .X(net1365),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1366 (.A(net1368),
    .X(net1366),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1367 (.A(net1368),
    .X(net1367),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1368 (.A(net1371),
    .X(net1368),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1370 (.A(net1371),
    .X(net1370),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1371 (.A(\i_ibex/id_stage_i/alu_op_b_mux_sel_dec ),
    .X(net1371),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1372 (.A(net1373),
    .X(net1372),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1373 (.A(\i_ibex/id_stage_i/alu_op_b_mux_sel_dec ),
    .X(net1373),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1374 (.A(net1376),
    .X(net1374),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1375 (.A(net1376),
    .X(net1375),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1376 (.A(\i_ibex/id_stage_i/alu_op_b_mux_sel_dec ),
    .X(net1376),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1377 (.A(net1378),
    .X(net1377),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1378 (.A(\i_ibex/id_stage_i/_0359_ ),
    .X(net1378),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1379 (.A(net1381),
    .X(net1379),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1380 (.A(net1381),
    .X(net1380),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1381 (.A(\i_ibex/id_stage_i/_0359_ ),
    .X(net1381),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1382 (.A(net1383),
    .X(net1382),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1383 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0182_ ),
    .X(net1383),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1384 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0152_ ),
    .X(net1384),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1385 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0126_ ),
    .X(net1385),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1386 (.A(net1387),
    .X(net1386),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1387 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0098_ ),
    .X(net1387),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1388 (.A(net1390),
    .X(net1388),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1389 (.A(net1390),
    .X(net1389),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1390 (.X(net1390),
    .A(net1393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1391 (.X(net1391),
    .A(net1393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1392 (.A(net1393),
    .X(net1392),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1393 (.A(\i_ibex/rf_we_lsu ),
    .X(net1393),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1394 (.X(net1394),
    .A(\i_ibex/id_stage_i/controller_i/_080_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1395 (.A(net1396),
    .X(net1395),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1396 (.A(\i_ibex/id_stage_i/controller_i/_038_ ),
    .X(net1396),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1397 (.A(net1398),
    .X(net1397),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1398 (.A(\i_ibex/cs_registers_i/minstret_counter_i/_0097_ ),
    .X(net1398),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1399 (.A(\i_ibex/load_store_unit_i/_0326_ ),
    .X(net1399),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1400 (.A(net1401),
    .X(net1400),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1401 (.A(\i_ibex/load_store_unit_i/_0216_ ),
    .X(net1401),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1402 (.A(net1403),
    .X(net1402),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1403 (.A(\i_ibex/load_store_unit_i/_0216_ ),
    .X(net1403),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1404 (.X(net1404),
    .A(net1408),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1405 (.A(net1408),
    .X(net1405),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1406 (.X(net1406),
    .A(net1407),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1407 (.X(net1407),
    .A(net1408),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1408 (.A(\i_ibex/id_stage_i/controller_i/_045_ ),
    .X(net1408),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1409 (.A(net1411),
    .X(net1409),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1410 (.A(net1411),
    .X(net1410),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1411 (.A(\i_ibex/load_store_unit_i/_0222_ ),
    .X(net1411),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1412 (.A(\i_ibex/load_store_unit_i/_0222_ ),
    .X(net1412),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1413 (.A(\i_ibex/load_store_unit_i/_0222_ ),
    .X(net1413),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1414 (.A(net1415),
    .X(net1414),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1415 (.A(net1422),
    .X(net1415),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1416 (.A(net1422),
    .X(net1416),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1417 (.A(net1422),
    .X(net1417),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1418 (.A(net1421),
    .X(net1418),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1419 (.A(net1421),
    .X(net1419),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1420 (.A(net1421),
    .X(net1420),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1421 (.A(net1422),
    .X(net1421),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1422 (.A(\i_ibex/load_store_unit_i/_0219_ ),
    .X(net1422),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1423 (.A(net1427),
    .X(net1423),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1424 (.A(net1427),
    .X(net1424),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1425 (.A(net1427),
    .X(net1425),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1426 (.A(net1427),
    .X(net1426),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1427 (.A(\i_ibex/load_store_unit_i/_0211_ ),
    .X(net1427),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1428 (.A(net1431),
    .X(net1428),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1429 (.A(net1431),
    .X(net1429),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1430 (.A(net1431),
    .X(net1430),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1431 (.A(\i_ibex/load_store_unit_i/_0211_ ),
    .X(net1431),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1432 (.A(net1435),
    .X(net1432),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1433 (.A(net1434),
    .X(net1433),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1434 (.A(net1435),
    .X(net1434),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1435 (.A(net1437),
    .X(net1435),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1436 (.A(net1437),
    .X(net1436),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1437 (.A(\i_ibex/load_store_unit_i/_0208_ ),
    .X(net1437),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1438 (.X(net1438),
    .A(net1439),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1439 (.X(net1439),
    .A(net1442),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1440 (.X(net1440),
    .A(net1441),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1441 (.X(net1441),
    .A(net1442),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1442 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_165_ ),
    .X(net1442),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1443 (.A(net1444),
    .X(net1443),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1444 (.A(net1447),
    .X(net1444),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1445 (.X(net1445),
    .A(net1447),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1446 (.X(net1446),
    .A(net1447),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1447 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_146_ ),
    .X(net1447),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1448 (.A(\i_ibex/id_stage_i/controller_i/_117_ ),
    .X(net1448),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1449 (.A(\i_ibex/id_stage_i/controller_i/_117_ ),
    .X(net1449),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1450 (.A(net1452),
    .X(net1450),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1451 (.A(net1452),
    .X(net1451),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1452 (.A(\i_ibex/id_stage_i/controller_i/_008_ ),
    .X(net1452),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1453 (.A(net1455),
    .X(net1453),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1454 (.A(net1455),
    .X(net1454),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1455 (.A(\i_ibex/id_stage_i/controller_i/_008_ ),
    .X(net1455),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1456 (.X(net1456),
    .A(\i_ibex/load_store_unit_i/_0242_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1457 (.A(\i_ibex/load_store_unit_i/_0235_ ),
    .X(net1457),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1458 (.A(\i_ibex/load_store_unit_i/rdata_offset_q_$_NOT__A_1_Y ),
    .X(net1458),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1459 (.A(\i_ibex/load_store_unit_i/ls_fsm_cs [2]),
    .X(net1459),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1460 (.A(\i_ibex/load_store_unit_i/ls_fsm_cs [1]),
    .X(net1460),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1461 (.A(\i_ibex/load_store_unit_i/ls_fsm_cs [1]),
    .X(net1461),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1462 (.A(\i_ibex/load_store_unit_i/ls_fsm_cs [0]),
    .X(net1462),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1463 (.A(\i_ibex/load_store_unit_i/ls_fsm_cs [0]),
    .X(net1463),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1464 (.A(\i_ibex/load_store_unit_i/handle_misaligned_q ),
    .X(net1464),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1465 (.X(net1465),
    .A(net1466),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1466 (.X(net1466),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/valid_req_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1467 (.X(net1467),
    .A(net1469),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1468 (.A(net1469),
    .X(net1468),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1469 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/valid_req_q ),
    .X(net1469),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1470 (.A(net1472),
    .X(net1470),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1471 (.A(net1472),
    .X(net1471),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1472 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_q [0]),
    .X(net1472),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1473 (.X(net1473),
    .A(net1476),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1474 (.X(net1474),
    .A(net1475),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1475 (.A(net1476),
    .X(net1475),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1476 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/valid_q [0]),
    .X(net1476),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1477 (.X(net1477),
    .A(net1478),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1478 (.X(net1478),
    .A(\i_ibex/pc_if [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1479 (.X(net1479),
    .A(net1484),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1480 (.A(net1484),
    .X(net1480),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1481 (.X(net1481),
    .A(net1483),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1482 (.X(net1482),
    .A(net1483),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1483 (.X(net1483),
    .A(net1484),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1484 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_busy [1]),
    .X(net1484),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1485 (.X(net1485),
    .A(\i_ibex/id_stage_i/controller_i/illegal_insn_q ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1486 (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [2]),
    .X(net1486),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1487 (.A(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A ),
    .X(net1487),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1488 (.A(\i_ibex/id_stage_i/controller_i/debug_single_step_i_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A ),
    .X(net1488),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1489 (.A(net1490),
    .X(net1489),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1490 (.A(\i_ibex/id_stage_i/controller_i/ctrl_fsm_cs [0]),
    .X(net1490),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1491 (.A(\i_ibex/cs_registers_i/minstret_raw [20]),
    .X(net1491),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1492 (.A(\i_ibex/cs_registers_i/minstret_raw [17]),
    .X(net1492),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1493 (.A(net1494),
    .X(net1493),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1494 (.A(\i_ibex/cs_registers_i/minstret_raw [16]),
    .X(net1494),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1495 (.X(net1495),
    .A(net1496),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1496 (.X(net1496),
    .A(\i_ibex/ex_block_i/alu_i/_0706_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 load_slew1497 (.X(net1497),
    .A(net1637),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 load_slew1498 (.X(net1498),
    .A(net1637),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 load_slew1499 (.X(net1499),
    .A(net1554),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 load_slew1500 (.X(net1500),
    .A(net1640),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 load_slew1501 (.A(rst_ni),
    .X(net1501),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 load_slew1502 (.X(net1502),
    .A(rst_ni),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1503 (.X(net1503),
    .A(net1504),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1504 (.X(net1504),
    .A(net1507),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1505 (.X(net1505),
    .A(net1507),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1506 (.X(net1506),
    .A(net1507),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1507 (.A(net282),
    .X(net1507),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1508 (.X(net1508),
    .A(net1512),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1509 (.X(net1509),
    .A(net1512),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1510 (.X(net1510),
    .A(net1512),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1511 (.X(net1511),
    .A(net1512),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout1512 (.A(net256),
    .X(net1512),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1513 (.A(\i_ibex/rf_rdata_b [0]),
    .X(net1513),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1514 (.A(\i_ibex/alu_operand_a_ex [0]),
    .X(net1514),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 rebuffer1515 (.X(net1515),
    .A(\i_ibex/cs_registers_i/mcycle_counter_i/_216_ ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1516 (.A(\i_ibex/ex_block_i/alu_i/_0899_ ),
    .X(net1516),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_regs_0_clk_sys (.A(clk_i),
    .X(delaynet_0_clk_sys),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_0_clk_i_regs (.X(clknet_leaf_0_clk_i_regs),
    .A(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_1_clk_i_regs (.X(clknet_leaf_1_clk_i_regs),
    .A(clknet_5_2__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_2_clk_i_regs (.X(clknet_leaf_2_clk_i_regs),
    .A(clknet_5_3__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_3_clk_i_regs (.X(clknet_leaf_3_clk_i_regs),
    .A(clknet_5_2__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_4_clk_i_regs (.X(clknet_leaf_4_clk_i_regs),
    .A(clknet_5_3__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_5_clk_i_regs (.X(clknet_leaf_5_clk_i_regs),
    .A(clknet_5_3__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_6_clk_i_regs (.X(clknet_leaf_6_clk_i_regs),
    .A(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_7_clk_i_regs (.X(clknet_leaf_7_clk_i_regs),
    .A(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_8_clk_i_regs (.X(clknet_leaf_8_clk_i_regs),
    .A(clknet_5_2__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_9_clk_i_regs (.X(clknet_leaf_9_clk_i_regs),
    .A(clknet_5_2__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_10_clk_i_regs (.X(clknet_leaf_10_clk_i_regs),
    .A(clknet_5_2__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_11_clk_i_regs (.X(clknet_leaf_11_clk_i_regs),
    .A(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_12_clk_i_regs (.X(clknet_leaf_12_clk_i_regs),
    .A(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_13_clk_i_regs (.X(clknet_leaf_13_clk_i_regs),
    .A(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_14_clk_i_regs (.X(clknet_leaf_14_clk_i_regs),
    .A(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_15_clk_i_regs (.X(clknet_leaf_15_clk_i_regs),
    .A(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_16_clk_i_regs (.X(clknet_leaf_16_clk_i_regs),
    .A(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_17_clk_i_regs (.X(clknet_leaf_17_clk_i_regs),
    .A(clknet_5_10__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_18_clk_i_regs (.X(clknet_leaf_18_clk_i_regs),
    .A(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_19_clk_i_regs (.X(clknet_leaf_19_clk_i_regs),
    .A(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_20_clk_i_regs (.X(clknet_leaf_20_clk_i_regs),
    .A(clknet_5_11__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_21_clk_i_regs (.X(clknet_leaf_21_clk_i_regs),
    .A(clknet_5_12__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_22_clk_i_regs (.X(clknet_leaf_22_clk_i_regs),
    .A(clknet_5_12__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_23_clk_i_regs (.X(clknet_leaf_23_clk_i_regs),
    .A(clknet_5_12__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_24_clk_i_regs (.X(clknet_leaf_24_clk_i_regs),
    .A(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_25_clk_i_regs (.X(clknet_leaf_25_clk_i_regs),
    .A(clknet_5_12__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_27_clk_i_regs (.X(clknet_leaf_27_clk_i_regs),
    .A(clknet_5_3__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_28_clk_i_regs (.X(clknet_leaf_28_clk_i_regs),
    .A(clknet_5_6__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_29_clk_i_regs (.X(clknet_leaf_29_clk_i_regs),
    .A(clknet_5_6__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_30_clk_i_regs (.X(clknet_leaf_30_clk_i_regs),
    .A(clknet_5_7__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_31_clk_i_regs (.X(clknet_leaf_31_clk_i_regs),
    .A(clknet_5_13__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_32_clk_i_regs (.X(clknet_leaf_32_clk_i_regs),
    .A(clknet_5_13__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_33_clk_i_regs (.X(clknet_leaf_33_clk_i_regs),
    .A(clknet_5_13__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_34_clk_i_regs (.X(clknet_leaf_34_clk_i_regs),
    .A(clknet_5_13__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_35_clk_i_regs (.X(clknet_leaf_35_clk_i_regs),
    .A(clknet_5_13__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_36_clk_i_regs (.X(clknet_leaf_36_clk_i_regs),
    .A(clknet_5_29__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_37_clk_i_regs (.X(clknet_leaf_37_clk_i_regs),
    .A(clknet_5_15__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_38_clk_i_regs (.X(clknet_leaf_38_clk_i_regs),
    .A(clknet_5_15__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_39_clk_i_regs (.X(clknet_leaf_39_clk_i_regs),
    .A(clknet_5_15__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_40_clk_i_regs (.X(clknet_leaf_40_clk_i_regs),
    .A(clknet_5_15__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_41_clk_i_regs (.X(clknet_leaf_41_clk_i_regs),
    .A(clknet_5_15__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_42_clk_i_regs (.X(clknet_leaf_42_clk_i_regs),
    .A(clknet_5_28__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_43_clk_i_regs (.X(clknet_leaf_43_clk_i_regs),
    .A(clknet_5_25__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_45_clk_i_regs (.X(clknet_leaf_45_clk_i_regs),
    .A(clknet_5_14__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_46_clk_i_regs (.X(clknet_leaf_46_clk_i_regs),
    .A(clknet_5_14__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_47_clk_i_regs (.X(clknet_leaf_47_clk_i_regs),
    .A(clknet_5_14__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_48_clk_i_regs (.X(clknet_leaf_48_clk_i_regs),
    .A(clknet_5_12__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_49_clk_i_regs (.X(clknet_leaf_49_clk_i_regs),
    .A(clknet_5_14__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_50_clk_i_regs (.X(clknet_leaf_50_clk_i_regs),
    .A(clknet_5_14__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_51_clk_i_regs (.X(clknet_leaf_51_clk_i_regs),
    .A(clknet_5_11__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_52_clk_i_regs (.X(clknet_leaf_52_clk_i_regs),
    .A(clknet_5_11__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_53_clk_i_regs (.X(clknet_leaf_53_clk_i_regs),
    .A(clknet_5_11__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_54_clk_i_regs (.X(clknet_leaf_54_clk_i_regs),
    .A(clknet_5_10__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_55_clk_i_regs (.X(clknet_leaf_55_clk_i_regs),
    .A(clknet_5_10__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_56_clk_i_regs (.X(clknet_leaf_56_clk_i_regs),
    .A(clknet_5_10__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_57_clk_i_regs (.X(clknet_leaf_57_clk_i_regs),
    .A(clknet_5_10__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_58_clk_i_regs (.X(clknet_leaf_58_clk_i_regs),
    .A(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_59_clk_i_regs (.X(clknet_leaf_59_clk_i_regs),
    .A(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_60_clk_i_regs (.X(clknet_leaf_60_clk_i_regs),
    .A(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_61_clk_i_regs (.X(clknet_leaf_61_clk_i_regs),
    .A(clknet_5_11__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_62_clk_i_regs (.X(clknet_leaf_62_clk_i_regs),
    .A(clknet_5_25__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_63_clk_i_regs (.X(clknet_leaf_63_clk_i_regs),
    .A(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_64_clk_i_regs (.X(clknet_leaf_64_clk_i_regs),
    .A(clknet_5_25__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_65_clk_i_regs (.X(clknet_leaf_65_clk_i_regs),
    .A(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_66_clk_i_regs (.X(clknet_leaf_66_clk_i_regs),
    .A(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_67_clk_i_regs (.X(clknet_leaf_67_clk_i_regs),
    .A(clknet_5_26__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_68_clk_i_regs (.X(clknet_leaf_68_clk_i_regs),
    .A(clknet_5_26__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_69_clk_i_regs (.X(clknet_leaf_69_clk_i_regs),
    .A(clknet_5_26__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_70_clk_i_regs (.X(clknet_leaf_70_clk_i_regs),
    .A(clknet_5_26__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_71_clk_i_regs (.X(clknet_leaf_71_clk_i_regs),
    .A(clknet_5_26__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_72_clk_i_regs (.X(clknet_leaf_72_clk_i_regs),
    .A(clknet_5_27__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_73_clk_i_regs (.X(clknet_leaf_73_clk_i_regs),
    .A(clknet_5_27__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_74_clk_i_regs (.X(clknet_leaf_74_clk_i_regs),
    .A(clknet_5_27__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_75_clk_i_regs (.X(clknet_leaf_75_clk_i_regs),
    .A(clknet_5_30__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_76_clk_i_regs (.X(clknet_leaf_76_clk_i_regs),
    .A(clknet_5_27__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_77_clk_i_regs (.X(clknet_leaf_77_clk_i_regs),
    .A(clknet_5_27__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_78_clk_i_regs (.X(clknet_leaf_78_clk_i_regs),
    .A(clknet_5_30__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_79_clk_i_regs (.X(clknet_leaf_79_clk_i_regs),
    .A(clknet_5_25__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_80_clk_i_regs (.X(clknet_leaf_80_clk_i_regs),
    .A(clknet_5_28__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_81_clk_i_regs (.X(clknet_leaf_81_clk_i_regs),
    .A(clknet_5_30__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_82_clk_i_regs (.X(clknet_leaf_82_clk_i_regs),
    .A(clknet_5_28__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_83_clk_i_regs (.X(clknet_leaf_83_clk_i_regs),
    .A(clknet_5_31__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_84_clk_i_regs (.X(clknet_leaf_84_clk_i_regs),
    .A(clknet_5_30__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_85_clk_i_regs (.X(clknet_leaf_85_clk_i_regs),
    .A(clknet_5_30__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_86_clk_i_regs (.X(clknet_leaf_86_clk_i_regs),
    .A(clknet_5_31__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_87_clk_i_regs (.X(clknet_leaf_87_clk_i_regs),
    .A(clknet_5_31__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_88_clk_i_regs (.X(clknet_leaf_88_clk_i_regs),
    .A(clknet_5_31__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_89_clk_i_regs (.X(clknet_leaf_89_clk_i_regs),
    .A(clknet_5_31__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_91_clk_i_regs (.X(clknet_leaf_91_clk_i_regs),
    .A(clknet_5_16__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_92_clk_i_regs (.X(clknet_leaf_92_clk_i_regs),
    .A(clknet_5_29__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_93_clk_i_regs (.X(clknet_leaf_93_clk_i_regs),
    .A(clknet_5_28__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_94_clk_i_regs (.X(clknet_leaf_94_clk_i_regs),
    .A(clknet_5_28__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_95_clk_i_regs (.X(clknet_leaf_95_clk_i_regs),
    .A(clknet_5_29__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_96_clk_i_regs (.X(clknet_leaf_96_clk_i_regs),
    .A(clknet_5_29__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_97_clk_i_regs (.X(clknet_leaf_97_clk_i_regs),
    .A(clknet_5_16__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_98_clk_i_regs (.X(clknet_leaf_98_clk_i_regs),
    .A(clknet_5_16__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_99_clk_i_regs (.X(clknet_leaf_99_clk_i_regs),
    .A(clknet_5_16__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_103_clk_i_regs (.X(clknet_leaf_103_clk_i_regs),
    .A(clknet_5_18__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_104_clk_i_regs (.X(clknet_leaf_104_clk_i_regs),
    .A(clknet_5_18__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_105_clk_i_regs (.X(clknet_leaf_105_clk_i_regs),
    .A(clknet_5_18__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_106_clk_i_regs (.X(clknet_leaf_106_clk_i_regs),
    .A(clknet_5_19__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_107_clk_i_regs (.X(clknet_leaf_107_clk_i_regs),
    .A(clknet_5_19__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_108_clk_i_regs (.X(clknet_leaf_108_clk_i_regs),
    .A(clknet_5_19__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_109_clk_i_regs (.X(clknet_leaf_109_clk_i_regs),
    .A(clknet_5_19__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_110_clk_i_regs (.X(clknet_leaf_110_clk_i_regs),
    .A(clknet_5_19__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_111_clk_i_regs (.X(clknet_leaf_111_clk_i_regs),
    .A(clknet_5_18__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_112_clk_i_regs (.X(clknet_leaf_112_clk_i_regs),
    .A(clknet_5_18__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_113_clk_i_regs (.X(clknet_leaf_113_clk_i_regs),
    .A(clknet_5_22__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_114_clk_i_regs (.X(clknet_leaf_114_clk_i_regs),
    .A(clknet_5_22__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_115_clk_i_regs (.X(clknet_leaf_115_clk_i_regs),
    .A(clknet_5_22__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_116_clk_i_regs (.X(clknet_leaf_116_clk_i_regs),
    .A(clknet_5_22__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_117_clk_i_regs (.X(clknet_leaf_117_clk_i_regs),
    .A(clknet_5_22__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_118_clk_i_regs (.X(clknet_leaf_118_clk_i_regs),
    .A(clknet_5_23__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_119_clk_i_regs (.X(clknet_leaf_119_clk_i_regs),
    .A(clknet_5_23__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_120_clk_i_regs (.X(clknet_leaf_120_clk_i_regs),
    .A(clknet_5_23__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_121_clk_i_regs (.X(clknet_leaf_121_clk_i_regs),
    .A(clknet_5_23__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_122_clk_i_regs (.X(clknet_leaf_122_clk_i_regs),
    .A(clknet_5_23__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_123_clk_i_regs (.X(clknet_leaf_123_clk_i_regs),
    .A(clknet_5_21__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_124_clk_i_regs (.X(clknet_leaf_124_clk_i_regs),
    .A(clknet_5_21__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_125_clk_i_regs (.X(clknet_leaf_125_clk_i_regs),
    .A(clknet_5_21__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_126_clk_i_regs (.X(clknet_leaf_126_clk_i_regs),
    .A(clknet_5_21__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_128_clk_i_regs (.X(clknet_leaf_128_clk_i_regs),
    .A(clknet_5_17__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_129_clk_i_regs (.X(clknet_leaf_129_clk_i_regs),
    .A(clknet_5_17__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_130_clk_i_regs (.X(clknet_leaf_130_clk_i_regs),
    .A(clknet_5_20__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_131_clk_i_regs (.X(clknet_leaf_131_clk_i_regs),
    .A(clknet_5_21__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_132_clk_i_regs (.X(clknet_leaf_132_clk_i_regs),
    .A(clknet_5_20__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_133_clk_i_regs (.X(clknet_leaf_133_clk_i_regs),
    .A(clknet_5_20__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_134_clk_i_regs (.X(clknet_leaf_134_clk_i_regs),
    .A(clknet_5_20__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_135_clk_i_regs (.X(clknet_leaf_135_clk_i_regs),
    .A(clknet_5_17__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_137_clk_i_regs (.X(clknet_leaf_137_clk_i_regs),
    .A(clknet_5_7__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_138_clk_i_regs (.X(clknet_leaf_138_clk_i_regs),
    .A(clknet_5_7__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_139_clk_i_regs (.X(clknet_leaf_139_clk_i_regs),
    .A(clknet_5_6__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_140_clk_i_regs (.X(clknet_leaf_140_clk_i_regs),
    .A(clknet_5_6__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_141_clk_i_regs (.X(clknet_leaf_141_clk_i_regs),
    .A(clknet_5_7__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_142_clk_i_regs (.X(clknet_leaf_142_clk_i_regs),
    .A(clknet_5_7__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_143_clk_i_regs (.X(clknet_leaf_143_clk_i_regs),
    .A(clknet_5_5__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_144_clk_i_regs (.X(clknet_leaf_144_clk_i_regs),
    .A(clknet_5_5__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_145_clk_i_regs (.X(clknet_leaf_145_clk_i_regs),
    .A(clknet_5_5__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_146_clk_i_regs (.X(clknet_leaf_146_clk_i_regs),
    .A(clknet_5_4__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_147_clk_i_regs (.X(clknet_leaf_147_clk_i_regs),
    .A(clknet_5_4__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_148_clk_i_regs (.X(clknet_leaf_148_clk_i_regs),
    .A(clknet_5_5__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_149_clk_i_regs (.X(clknet_leaf_149_clk_i_regs),
    .A(clknet_5_5__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_150_clk_i_regs (.X(clknet_leaf_150_clk_i_regs),
    .A(clknet_5_4__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_151_clk_i_regs (.X(clknet_leaf_151_clk_i_regs),
    .A(clknet_5_6__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_152_clk_i_regs (.X(clknet_leaf_152_clk_i_regs),
    .A(clknet_5_4__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_153_clk_i_regs (.X(clknet_leaf_153_clk_i_regs),
    .A(clknet_5_4__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_154_clk_i_regs (.X(clknet_leaf_154_clk_i_regs),
    .A(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_155_clk_i_regs (.X(clknet_leaf_155_clk_i_regs),
    .A(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_156_clk_i_regs (.X(clknet_leaf_156_clk_i_regs),
    .A(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_157_clk_i_regs (.X(clknet_leaf_157_clk_i_regs),
    .A(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_158_clk_i_regs (.X(clknet_leaf_158_clk_i_regs),
    .A(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_159_clk_i_regs (.X(clknet_leaf_159_clk_i_regs),
    .A(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_160_clk_i_regs (.X(clknet_leaf_160_clk_i_regs),
    .A(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_161_clk_i_regs (.X(clknet_leaf_161_clk_i_regs),
    .A(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_162_clk_i_regs (.X(clknet_leaf_162_clk_i_regs),
    .A(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_163_clk_i_regs (.X(clknet_leaf_163_clk_i_regs),
    .A(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .X(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_0_0_clk_i_regs (.X(clknet_4_0_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_1_0_clk_i_regs (.X(clknet_4_1_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_2_0_clk_i_regs (.X(clknet_4_2_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_3_0_clk_i_regs (.X(clknet_4_3_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_4_0_clk_i_regs (.X(clknet_4_4_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_5_0_clk_i_regs (.X(clknet_4_5_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_6_0_clk_i_regs (.X(clknet_4_6_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_7_0_clk_i_regs (.X(clknet_4_7_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_8_0_clk_i_regs (.X(clknet_4_8_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_9_0_clk_i_regs (.X(clknet_4_9_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_10_0_clk_i_regs (.X(clknet_4_10_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_11_0_clk_i_regs (.X(clknet_4_11_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_12_0_clk_i_regs (.X(clknet_4_12_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_13_0_clk_i_regs (.X(clknet_4_13_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_14_0_clk_i_regs (.X(clknet_4_14_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_15_0_clk_i_regs (.X(clknet_4_15_0_clk_i_regs),
    .A(clknet_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_0__f_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .X(clknet_5_0__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_1__f_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .X(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_2__f_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .X(clknet_5_2__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_3__f_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .X(clknet_5_3__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_4__f_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .X(clknet_5_4__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_5__f_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .X(clknet_5_5__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_6__f_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .X(clknet_5_6__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_7__f_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .X(clknet_5_7__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_8__f_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .X(clknet_5_8__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_9__f_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .X(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_10__f_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .X(clknet_5_10__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_11__f_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .X(clknet_5_11__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_12__f_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .X(clknet_5_12__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_13__f_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .X(clknet_5_13__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_14__f_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .X(clknet_5_14__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_15__f_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .X(clknet_5_15__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_16__f_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .X(clknet_5_16__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_17__f_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .X(clknet_5_17__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_18__f_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .X(clknet_5_18__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_19__f_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .X(clknet_5_19__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_20__f_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .X(clknet_5_20__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_21__f_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .X(clknet_5_21__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_22__f_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .X(clknet_5_22__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_23__f_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .X(clknet_5_23__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_24__f_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .X(clknet_5_24__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_25__f_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .X(clknet_5_25__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_26__f_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .X(clknet_5_26__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_27__f_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .X(clknet_5_27__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_28__f_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .X(clknet_5_28__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_29__f_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .X(clknet_5_29__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_30__f_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .X(clknet_5_30__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_31__f_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .X(clknet_5_31__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload0 (.A(clknet_5_1__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload1 (.A(clknet_5_3__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload2 (.A(clknet_5_9__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload3 (.A(clknet_5_17__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload4 (.A(clknet_5_20__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_8 clkload5 (.A(clknet_5_25__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload6 (.A(clknet_5_29__leaf_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_0_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload8 (.VDD(VDD),
    .A(clknet_leaf_159_clk_i_regs),
    .VSS(VSS));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_160_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload10 (.VDD(VDD),
    .A(clknet_leaf_154_clk_i_regs),
    .VSS(VSS));
 sg13g2_buf_2 clkload11 (.A(clknet_leaf_155_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload12 (.A(clknet_leaf_157_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload13 (.A(clknet_leaf_158_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_1_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload15 (.A(clknet_leaf_3_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload16 (.A(clknet_leaf_9_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_10_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload18 (.A(clknet_leaf_2_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_4_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_27_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload21 (.A(clknet_leaf_146_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload22 (.A(clknet_leaf_147_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_150_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_152_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_143_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload26 (.A(clknet_leaf_144_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_148_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload28 (.A(clknet_leaf_149_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_28_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload30 (.A(clknet_leaf_29_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload31 (.A(clknet_leaf_140_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_151_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload33 (.A(clknet_leaf_30_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload34 (.A(clknet_leaf_137_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_138_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload36 (.A(clknet_leaf_142_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload37 (.A(clknet_leaf_11_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload38 (.A(clknet_leaf_13_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload39 (.A(clknet_leaf_14_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload40 (.A(clknet_leaf_15_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_16_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload42 (.VDD(VDD),
    .A(clknet_leaf_6_clk_i_regs),
    .VSS(VSS));
 sg13g2_buf_2 clkload43 (.A(clknet_leaf_7_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload44 (.A(clknet_leaf_19_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload45 (.A(clknet_leaf_24_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload46 (.A(clknet_leaf_54_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload47 (.A(clknet_leaf_55_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload48 (.A(clknet_leaf_56_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload49 (.VDD(VDD),
    .A(clknet_leaf_57_clk_i_regs),
    .VSS(VSS));
 sg13g2_buf_2 clkload50 (.A(clknet_leaf_20_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload51 (.A(clknet_leaf_51_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload52 (.A(clknet_leaf_52_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 clkload53 (.A(clknet_leaf_61_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload54 (.A(clknet_leaf_21_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload55 (.A(clknet_leaf_23_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload56 (.A(clknet_leaf_25_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload57 (.A(clknet_leaf_48_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload58 (.A(clknet_leaf_31_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload59 (.A(clknet_leaf_32_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 clkload60 (.A(clknet_leaf_33_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload61 (.A(clknet_leaf_35_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload62 (.A(clknet_leaf_46_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload63 (.A(clknet_leaf_47_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload64 (.A(clknet_leaf_49_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload65 (.VDD(VDD),
    .A(clknet_leaf_50_clk_i_regs),
    .VSS(VSS));
 sg13g2_inv_4 clkload66 (.A(clknet_leaf_38_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload67 (.A(clknet_leaf_39_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload68 (.A(clknet_leaf_40_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload69 (.A(clknet_leaf_41_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload70 (.A(clknet_leaf_91_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload71 (.A(clknet_leaf_97_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload72 (.A(clknet_leaf_98_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload73 (.A(clknet_leaf_128_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload74 (.A(clknet_leaf_135_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload75 (.A(clknet_leaf_103_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload76 (.A(clknet_leaf_104_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload77 (.A(clknet_leaf_105_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload78 (.A(clknet_leaf_111_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload79 (.A(clknet_leaf_106_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload80 (.A(clknet_leaf_108_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload81 (.A(clknet_leaf_109_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload82 (.A(clknet_leaf_110_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload83 (.A(clknet_leaf_132_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload84 (.A(clknet_leaf_133_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload85 (.A(clknet_leaf_134_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload86 (.A(clknet_leaf_125_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload87 (.A(clknet_leaf_126_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload88 (.A(clknet_leaf_131_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload89 (.A(clknet_leaf_114_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload90 (.A(clknet_leaf_115_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload91 (.A(clknet_leaf_116_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload92 (.A(clknet_leaf_117_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload93 (.A(clknet_leaf_118_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload94 (.A(clknet_leaf_120_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload95 (.VDD(VDD),
    .A(clknet_leaf_122_clk_i_regs),
    .VSS(VSS));
 sg13g2_inv_4 clkload96 (.A(clknet_leaf_59_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload97 (.A(clknet_leaf_60_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload98 (.A(clknet_leaf_63_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload99 (.A(clknet_leaf_65_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload100 (.VDD(VDD),
    .A(clknet_leaf_66_clk_i_regs),
    .VSS(VSS));
 sg13g2_inv_4 clkload101 (.A(clknet_leaf_62_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload102 (.A(clknet_leaf_64_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload103 (.A(clknet_leaf_79_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload104 (.A(clknet_leaf_67_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload105 (.A(clknet_leaf_69_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload106 (.A(clknet_leaf_71_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload107 (.A(clknet_leaf_72_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload108 (.A(clknet_leaf_73_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload109 (.A(clknet_leaf_76_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload110 (.A(clknet_leaf_77_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload111 (.A(clknet_leaf_42_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload112 (.A(clknet_leaf_80_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload113 (.A(clknet_leaf_82_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload114 (.A(clknet_leaf_93_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload115 (.A(clknet_leaf_36_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload116 (.A(clknet_leaf_92_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload117 (.A(clknet_leaf_96_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload118 (.A(clknet_leaf_78_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload119 (.VDD(VDD),
    .A(clknet_leaf_81_clk_i_regs),
    .VSS(VSS));
 sg13g2_buf_2 clkload120 (.A(clknet_leaf_84_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload121 (.A(clknet_leaf_83_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload122 (.A(clknet_leaf_86_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload123 (.A(clknet_leaf_87_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload124 (.A(clknet_leaf_88_clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 delaybuf_0_clk_sys (.A(delaynet_0_clk_sys),
    .X(delaynet_1_clk_sys),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 delaybuf_1_clk_sys (.A(delaynet_1_clk_sys),
    .X(delaynet_2_clk_sys),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 delaybuf_2_clk_sys (.A(delaynet_2_clk_sys),
    .X(clk_i_regs),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 rebuffer1517 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_155_ ),
    .X(net1517),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1518 (.A(\i_ibex/ex_block_i/alu_adder_result_ext [30]),
    .X(net1518),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1519 (.A(\i_ibex/ex_block_i/alu_adder_result_ext [29]),
    .X(net1519),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1520 (.A(\i_ibex/ex_block_i/alu_adder_result_ext [31]),
    .X(net1520),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 rebuffer1521 (.A(\i_ibex/ex_block_i/alu_i/_1176_ ),
    .X(net1521),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd1_1 rebuffer1522 (.A(net1521),
    .X(net1522),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1523 (.A(net1524),
    .X(net1523),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1524 (.A(net1525),
    .X(net1524),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1525 (.A(net1553),
    .X(net1525),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1526 (.A(net1527),
    .X(net1526),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1527 (.A(net1553),
    .X(net1527),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1528 (.A(net1529),
    .X(net1528),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1529 (.A(net1530),
    .X(net1529),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1530 (.A(net1552),
    .X(net1530),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1531 (.A(net1532),
    .X(net1531),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1532 (.A(net1533),
    .X(net1532),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1533 (.A(net1552),
    .X(net1533),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1534 (.A(net1536),
    .X(net1534),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1535 (.A(net1536),
    .X(net1535),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1536 (.A(net1551),
    .X(net1536),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1537 (.A(net1538),
    .X(net1537),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1538 (.A(net1539),
    .X(net1538),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1539 (.A(net1551),
    .X(net1539),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1540 (.A(net1544),
    .X(net1540),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1541 (.A(net1542),
    .X(net1541),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1542 (.A(net1544),
    .X(net1542),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1543 (.A(net1544),
    .X(net1543),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1544 (.A(net1551),
    .X(net1544),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1545 (.A(net1546),
    .X(net1545),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1546 (.A(net1550),
    .X(net1546),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1547 (.A(net1549),
    .X(net1547),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1548 (.A(net1549),
    .X(net1548),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1549 (.A(net1550),
    .X(net1549),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1550 (.A(net1551),
    .X(net1550),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1551 (.A(net1552),
    .X(net1551),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1552 (.A(net1553),
    .X(net1552),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1553 (.A(net1499),
    .X(net1553),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1554 (.A(net1556),
    .X(net1554),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1555 (.A(net1556),
    .X(net1555),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1556 (.A(net1557),
    .X(net1556),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1557 (.A(net1561),
    .X(net1557),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1558 (.A(net1559),
    .X(net1558),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1559 (.A(net1560),
    .X(net1559),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1560 (.A(net1561),
    .X(net1560),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1561 (.A(net1562),
    .X(net1561),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1562 (.A(net1500),
    .X(net1562),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1563 (.A(net1565),
    .X(net1563),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1564 (.A(net1565),
    .X(net1564),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1565 (.A(net1566),
    .X(net1565),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1566 (.A(net1567),
    .X(net1566),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1567 (.A(net1579),
    .X(net1567),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1568 (.A(net1570),
    .X(net1568),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1569 (.A(net1570),
    .X(net1569),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1570 (.A(net1579),
    .X(net1570),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1571 (.A(net1572),
    .X(net1571),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1572 (.A(net1574),
    .X(net1572),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1573 (.A(net1574),
    .X(net1573),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1574 (.A(net1579),
    .X(net1574),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1575 (.A(net1578),
    .X(net1575),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1576 (.A(net1578),
    .X(net1576),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1577 (.A(net1578),
    .X(net1577),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1578 (.A(net1579),
    .X(net1578),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1579 (.A(net1581),
    .X(net1579),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1580 (.A(net1581),
    .X(net1580),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1581 (.A(net1500),
    .X(net1581),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1582 (.A(net1583),
    .X(net1582),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1583 (.A(net1584),
    .X(net1583),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1584 (.A(net1613),
    .X(net1584),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1585 (.A(net1587),
    .X(net1585),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1586 (.A(net1587),
    .X(net1586),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1587 (.A(net1597),
    .X(net1587),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1588 (.A(net1591),
    .X(net1588),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1589 (.A(net1590),
    .X(net1589),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1590 (.A(net1591),
    .X(net1590),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1591 (.A(net1597),
    .X(net1591),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1592 (.A(net1594),
    .X(net1592),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1593 (.A(net1594),
    .X(net1593),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1594 (.A(net1595),
    .X(net1594),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1595 (.A(net1596),
    .X(net1595),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1596 (.A(net1597),
    .X(net1596),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1597 (.A(net1613),
    .X(net1597),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1598 (.A(net1601),
    .X(net1598),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1599 (.A(net1600),
    .X(net1599),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1600 (.A(net1601),
    .X(net1600),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1601 (.A(net1607),
    .X(net1601),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1602 (.A(net1607),
    .X(net1602),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1603 (.A(net1607),
    .X(net1603),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1604 (.A(net1605),
    .X(net1604),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1605 (.A(net1606),
    .X(net1605),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1606 (.A(net1607),
    .X(net1606),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1607 (.A(net1613),
    .X(net1607),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1608 (.A(net1612),
    .X(net1608),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1609 (.A(net1612),
    .X(net1609),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1610 (.A(net1612),
    .X(net1610),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1611 (.A(net1612),
    .X(net1611),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1612 (.A(net1613),
    .X(net1612),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1613 (.A(net1498),
    .X(net1613),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1614 (.A(net1615),
    .X(net1614),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1615 (.A(net1624),
    .X(net1615),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1616 (.A(net1618),
    .X(net1616),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1617 (.A(net1618),
    .X(net1617),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1618 (.A(net1624),
    .X(net1618),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1619 (.A(net1620),
    .X(net1619),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1620 (.A(net1622),
    .X(net1620),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1621 (.A(net1622),
    .X(net1621),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1622 (.A(net1624),
    .X(net1622),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1623 (.A(net1624),
    .X(net1623),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1624 (.A(net1636),
    .X(net1624),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1625 (.A(net1628),
    .X(net1625),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1626 (.A(net1628),
    .X(net1626),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1627 (.A(net1628),
    .X(net1627),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1628 (.A(net1636),
    .X(net1628),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1629 (.A(net1632),
    .X(net1629),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1630 (.A(net1632),
    .X(net1630),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1631 (.A(net1632),
    .X(net1631),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1632 (.A(net1635),
    .X(net1632),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1633 (.A(net1634),
    .X(net1633),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1634 (.A(net1635),
    .X(net1634),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1635 (.A(net1636),
    .X(net1635),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1636 (.A(net1497),
    .X(net1636),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1637 (.A(net1641),
    .X(net1637),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1638 (.A(net1640),
    .X(net1638),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1639 (.A(net1640),
    .X(net1639),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1640 (.A(net1641),
    .X(net1640),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1641 (.A(net1647),
    .X(net1641),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1642 (.A(net1643),
    .X(net1642),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1643 (.A(net1644),
    .X(net1643),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1644 (.A(net1647),
    .X(net1644),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1645 (.A(net1646),
    .X(net1645),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1646 (.A(net1647),
    .X(net1646),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1647 (.A(net1650),
    .X(net1647),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1648 (.A(net1650),
    .X(net1648),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1649 (.A(net1650),
    .X(net1649),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1650 (.A(net1656),
    .X(net1650),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1651 (.A(net1652),
    .X(net1651),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1652 (.A(net1653),
    .X(net1652),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1653 (.A(net1656),
    .X(net1653),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1654 (.A(net1655),
    .X(net1654),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1655 (.A(net1656),
    .X(net1655),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1656 (.A(net1502),
    .X(net1656),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1657 (.A(net1664),
    .X(net1657),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1658 (.A(net1659),
    .X(net1658),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1659 (.A(net1664),
    .X(net1659),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1660 (.A(net1661),
    .X(net1660),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1661 (.A(net1662),
    .X(net1661),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1662 (.A(net1663),
    .X(net1662),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1663 (.A(net1664),
    .X(net1663),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1664 (.A(net1502),
    .X(net1664),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1665 (.A(net1668),
    .X(net1665),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1666 (.A(net1667),
    .X(net1666),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1667 (.A(net1668),
    .X(net1667),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 fanout1668 (.A(net1670),
    .X(net1668),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 max_cap1669 (.X(net1669),
    .A(net1501),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_1 max_cap1670 (.A(net1501),
    .X(net1670),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd3_1 hold1671 (.A(instr_rvalid_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/branch_discard_s [1]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold1673 (.A(instr_gnt_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold1674 (.A(instr_rdata_i[28]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold1675 (.A(instr_rdata_i[3]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold1676 (.A(instr_rdata_i[17]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_113_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold1678 (.A(instr_rdata_i[18]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold1679 (.A(instr_rdata_i[4]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold1680 (.A(instr_rdata_i[22]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold1681 (.A(instr_rdata_i[15]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold1682 (.A(instr_rdata_i[21]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold1683 (.A(instr_rdata_i[25]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold1684 (.A(instr_rdata_i[14]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold1685 (.A(instr_rdata_i[29]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold1686 (.A(instr_rdata_i[23]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold1687 (.A(instr_rdata_i[11]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold1688 (.A(instr_rdata_i[8]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold1689 (.A(instr_rdata_i[6]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold1690 (.A(instr_rdata_i[19]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold1691 (.A(instr_rdata_i[1]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold1692 (.A(instr_rdata_i[26]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold1693 (.A(instr_rdata_i[24]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold1694 (.A(data_rdata_i[28]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\i_ibex/load_store_unit_i/_0056_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold1696 (.A(instr_rdata_i[7]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold1697 (.A(instr_rdata_i[20]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold1698 (.A(instr_rdata_i[0]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold1699 (.A(instr_err_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold1700 (.A(instr_rdata_i[27]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold1701 (.A(instr_rdata_i[31]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold1702 (.A(instr_rdata_i[12]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold1703 (.A(instr_rdata_i[30]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold1704 (.A(data_rdata_i[20]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\i_ibex/load_store_unit_i/_0047_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold1706 (.A(data_rdata_i[8]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\i_ibex/load_store_unit_i/_0044_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold1708 (.A(instr_rdata_i[13]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold1709 (.A(instr_rdata_i[16]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold1710 (.A(instr_rdata_i[10]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold1711 (.A(data_rdata_i[22]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\i_ibex/load_store_unit_i/_0049_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold1713 (.A(data_rdata_i[13]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\i_ibex/load_store_unit_i/_0063_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold1715 (.A(data_rdata_i[14]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\i_ibex/load_store_unit_i/_0064_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold1717 (.A(data_rdata_i[21]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\i_ibex/load_store_unit_i/_0048_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold1719 (.A(instr_rdata_i[2]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold1720 (.A(data_rdata_i[27]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\i_ibex/load_store_unit_i/_0054_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold1722 (.A(data_rdata_i[17]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\i_ibex/load_store_unit_i/_0067_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold1724 (.A(instr_rdata_i[9]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold1725 (.A(data_rdata_i[25]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\i_ibex/load_store_unit_i/_0052_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold1727 (.A(data_rdata_i[19]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\i_ibex/load_store_unit_i/_0046_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold1729 (.A(data_rdata_i[29]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\i_ibex/load_store_unit_i/_0057_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold1731 (.A(data_rdata_i[18]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\i_ibex/load_store_unit_i/_0045_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold1733 (.A(data_rdata_i[11]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\i_ibex/load_store_unit_i/_0061_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold1735 (.A(instr_rdata_i[5]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold1736 (.A(data_rdata_i[10]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\i_ibex/load_store_unit_i/_0060_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold1738 (.A(debug_req_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold1739 (.A(data_rdata_i[30]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\i_ibex/load_store_unit_i/_0058_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold1741 (.A(data_rdata_i[24]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold1742 (.A(data_rdata_i[12]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\i_ibex/load_store_unit_i/_0062_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold1744 (.A(data_rdata_i[31]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold1745 (.A(data_rdata_i[26]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold1746 (.A(data_rdata_i[9]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\i_ibex/load_store_unit_i/_0055_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold1748 (.A(data_rdata_i[16]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\i_ibex/load_store_unit_i/_0066_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold1750 (.A(data_rdata_i[23]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\i_ibex/load_store_unit_i/_0050_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold1752 (.A(data_rdata_i[15]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\i_ibex/load_store_unit_i/_0065_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold1754 (.A(data_gnt_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\i_ibex/load_store_unit_i/_0184_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\i_ibex/load_store_unit_i/_0037_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold1757 (.A(data_err_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\i_ibex/load_store_unit_i/_0040_ ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold1759 (.A(boot_addr_i[25]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold1760 (.A(boot_addr_i[18]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold1761 (.A(boot_addr_i[9]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold1762 (.A(boot_addr_i[20]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold1763 (.A(boot_addr_i[11]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold1764 (.A(boot_addr_i[12]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold1765 (.A(boot_addr_i[30]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold1766 (.A(boot_addr_i[24]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold1767 (.A(boot_addr_i[10]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold1768 (.A(boot_addr_i[23]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold1769 (.A(data_rvalid_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold1770 (.A(boot_addr_i[26]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold1771 (.A(boot_addr_i[31]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold1772 (.A(boot_addr_i[22]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold1773 (.A(boot_addr_i[17]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold1774 (.A(boot_addr_i[13]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold1775 (.A(boot_addr_i[21]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold1776 (.A(boot_addr_i[29]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold1777 (.A(boot_addr_i[28]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold1778 (.A(boot_addr_i[19]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold1779 (.A(boot_addr_i[8]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold1780 (.A(boot_addr_i[15]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold1781 (.A(boot_addr_i[27]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold1782 (.A(boot_addr_i[16]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold1783 (.A(boot_addr_i[14]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold1784 (.A(fetch_enable_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold1785 (.A(data_rvalid_i),
    .VDD(VDD),
    .VSS(VSS),
    .X(net1785));
 sg13g2_antennanp ANTENNA_1 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[11]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[13]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[15]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[16]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[17]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[18]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[19]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[20]));
 sg13g2_antennanp ANTENNA_18 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[21]));
 sg13g2_antennanp ANTENNA_19 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[22]));
 sg13g2_antennanp ANTENNA_20 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[23]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[25]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_25 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_26 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[27]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[28]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[29]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_30 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_31 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[31]));
 sg13g2_antennanp ANTENNA_32 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[9]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_34 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_35 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_36 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_37 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_38 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_39 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_40 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_41 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_42 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_43 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_44 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_45 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_46 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_47 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_48 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_49 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_50 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_51 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_52 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_53 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_54 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_55 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_56 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_57 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_58 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_59 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_60 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_61 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_62 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_63 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_64 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_65 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_66 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_67 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_68 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_69 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_70 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_71 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_72 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_73 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_74 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_75 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_76 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_77 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_78 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_79 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_80 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_81 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_82 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_83 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_84 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_85 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_86 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_87 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_88 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_89 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_90 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_91 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_92 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_93 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_94 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_95 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_96 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_97 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_98 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_99 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_100 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_101 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_102 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_103 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_104 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_105 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_106 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_107 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_108 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_109 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_110 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_111 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_112 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_113 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_114 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_115 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_116 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_117 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_118 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_119 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_120 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_121 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_122 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_123 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_124 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_125 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_126 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_127 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_128 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_129 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_130 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_131 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_132 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_133 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_134 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[10]));
 sg13g2_antennanp ANTENNA_135 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[11]));
 sg13g2_antennanp ANTENNA_136 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[12]));
 sg13g2_antennanp ANTENNA_137 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[13]));
 sg13g2_antennanp ANTENNA_138 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[14]));
 sg13g2_antennanp ANTENNA_139 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[15]));
 sg13g2_antennanp ANTENNA_140 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[16]));
 sg13g2_antennanp ANTENNA_141 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[17]));
 sg13g2_antennanp ANTENNA_142 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[17]));
 sg13g2_antennanp ANTENNA_143 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[18]));
 sg13g2_antennanp ANTENNA_144 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[19]));
 sg13g2_antennanp ANTENNA_145 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[20]));
 sg13g2_antennanp ANTENNA_146 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[21]));
 sg13g2_antennanp ANTENNA_147 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[22]));
 sg13g2_antennanp ANTENNA_148 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[23]));
 sg13g2_antennanp ANTENNA_149 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[24]));
 sg13g2_antennanp ANTENNA_150 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[25]));
 sg13g2_antennanp ANTENNA_151 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_152 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[27]));
 sg13g2_antennanp ANTENNA_153 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[28]));
 sg13g2_antennanp ANTENNA_154 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[29]));
 sg13g2_antennanp ANTENNA_155 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[2]));
 sg13g2_antennanp ANTENNA_156 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_157 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[31]));
 sg13g2_antennanp ANTENNA_158 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[3]));
 sg13g2_antennanp ANTENNA_159 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[3]));
 sg13g2_antennanp ANTENNA_160 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[4]));
 sg13g2_antennanp ANTENNA_161 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[5]));
 sg13g2_antennanp ANTENNA_162 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[6]));
 sg13g2_antennanp ANTENNA_163 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[7]));
 sg13g2_antennanp ANTENNA_164 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[8]));
 sg13g2_antennanp ANTENNA_165 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[9]));
 sg13g2_antennanp ANTENNA_166 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_gnt_i));
 sg13g2_antennanp ANTENNA_167 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[13]));
 sg13g2_antennanp ANTENNA_168 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[13]));
 sg13g2_antennanp ANTENNA_169 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[19]));
 sg13g2_antennanp ANTENNA_170 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[19]));
 sg13g2_antennanp ANTENNA_171 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_172 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_173 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_174 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_175 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_176 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_177 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_178 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_179 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_180 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[2]));
 sg13g2_antennanp ANTENNA_181 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_182 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_183 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_184 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_185 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[9]));
 sg13g2_antennanp ANTENNA_186 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[9]));
 sg13g2_antennanp ANTENNA_187 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_188 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_189 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_190 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_191 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_192 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_193 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_194 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_195 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_196 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_197 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_198 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_199 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_200 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[3]));
 sg13g2_antennanp ANTENNA_201 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[3]));
 sg13g2_antennanp ANTENNA_202 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_busy ));
 sg13g2_antennanp ANTENNA_203 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_204 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_205 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_206 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_207 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/pc_mux_id [1]));
 sg13g2_antennanp ANTENNA_208 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/perf_instr_ret_wb ));
 sg13g2_antennanp ANTENNA_209 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_210 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_211 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_212 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_213 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_214 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_215 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_216 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_217 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_218 (.VDD(VDD),
    .VSS(VSS),
    .A(net946));
 sg13g2_antennanp ANTENNA_219 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_220 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_221 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [17]));
 sg13g2_antennanp ANTENNA_222 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [17]));
 sg13g2_antennanp ANTENNA_223 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [17]));
 sg13g2_antennanp ANTENNA_224 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [17]));
 sg13g2_antennanp ANTENNA_225 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [25]));
 sg13g2_antennanp ANTENNA_226 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [25]));
 sg13g2_antennanp ANTENNA_227 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/ex_block_i/alu_adder_result_ext [25]));
 sg13g2_antennanp ANTENNA_228 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/id_stage_i/_0455_ ));
 sg13g2_antennanp ANTENNA_229 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/id_stage_i/_0462_ ));
 sg13g2_antennanp ANTENNA_230 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_231 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_232 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_233 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_234 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_235 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_236 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_237 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_238 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_239 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_240 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_241 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_242 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_243 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_244 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_245 (.VDD(VDD),
    .VSS(VSS),
    .A(net1497));
 sg13g2_antennanp ANTENNA_246 (.VDD(VDD),
    .VSS(VSS),
    .A(net1497));
 sg13g2_antennanp ANTENNA_247 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_248 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_249 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_250 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_251 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_252 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_253 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_254 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_255 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_256 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_257 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_258 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_259 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_260 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_261 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_262 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_263 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_264 (.VDD(VDD),
    .VSS(VSS),
    .A(net1664));
 sg13g2_antennanp ANTENNA_265 (.VDD(VDD),
    .VSS(VSS),
    .A(net1664));
 sg13g2_antennanp ANTENNA_266 (.VDD(VDD),
    .VSS(VSS),
    .A(net1664));
 sg13g2_antennanp ANTENNA_267 (.VDD(VDD),
    .VSS(VSS),
    .A(net1664));
 sg13g2_antennanp ANTENNA_268 (.VDD(VDD),
    .VSS(VSS),
    .A(net1664));
 sg13g2_antennanp ANTENNA_269 (.VDD(VDD),
    .VSS(VSS),
    .A(net1664));
 sg13g2_antennanp ANTENNA_270 (.VDD(VDD),
    .VSS(VSS),
    .A(net1720));
 sg13g2_antennanp ANTENNA_271 (.VDD(VDD),
    .VSS(VSS),
    .A(net1736));
 sg13g2_antennanp ANTENNA_272 (.VDD(VDD),
    .VSS(VSS),
    .A(net1742));
 sg13g2_antennanp ANTENNA_273 (.VDD(VDD),
    .VSS(VSS),
    .A(net1752));
 sg13g2_antennanp ANTENNA_274 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 sg13g2_antennanp ANTENNA_275 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_276 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_277 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_278 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_279 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_280 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_281 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[11]));
 sg13g2_antennanp ANTENNA_282 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_283 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_284 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[13]));
 sg13g2_antennanp ANTENNA_285 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_286 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_287 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[15]));
 sg13g2_antennanp ANTENNA_288 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[16]));
 sg13g2_antennanp ANTENNA_289 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[17]));
 sg13g2_antennanp ANTENNA_290 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[18]));
 sg13g2_antennanp ANTENNA_291 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[19]));
 sg13g2_antennanp ANTENNA_292 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[20]));
 sg13g2_antennanp ANTENNA_293 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[21]));
 sg13g2_antennanp ANTENNA_294 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[23]));
 sg13g2_antennanp ANTENNA_295 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_296 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_297 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[25]));
 sg13g2_antennanp ANTENNA_298 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_299 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_300 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[27]));
 sg13g2_antennanp ANTENNA_301 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[28]));
 sg13g2_antennanp ANTENNA_302 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[29]));
 sg13g2_antennanp ANTENNA_303 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_304 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_305 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[31]));
 sg13g2_antennanp ANTENNA_306 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[9]));
 sg13g2_antennanp ANTENNA_307 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_308 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_309 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_310 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_311 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_312 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_313 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_314 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_315 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_316 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_317 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_318 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_319 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_320 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_321 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_322 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_323 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_324 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_325 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_326 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_327 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_328 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_329 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_330 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_331 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_332 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_333 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_334 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_335 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_336 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_337 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_338 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_339 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_340 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_341 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_342 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_343 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_344 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_345 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[18]));
 sg13g2_antennanp ANTENNA_346 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_347 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_348 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_349 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_350 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_351 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_352 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_353 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_354 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_355 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_356 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_357 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_358 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_359 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_360 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_361 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_362 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_363 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_364 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_365 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_366 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_367 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[24]));
 sg13g2_antennanp ANTENNA_368 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[24]));
 sg13g2_antennanp ANTENNA_369 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[24]));
 sg13g2_antennanp ANTENNA_370 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[24]));
 sg13g2_antennanp ANTENNA_371 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_372 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_373 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_374 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_375 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_376 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_377 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_378 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_379 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[26]));
 sg13g2_antennanp ANTENNA_380 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_381 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_382 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_383 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_384 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_385 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_386 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_387 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_388 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_389 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[29]));
 sg13g2_antennanp ANTENNA_390 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_391 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_392 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_393 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_394 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_395 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_396 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_397 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_398 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_399 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_400 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_401 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_402 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_403 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_404 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_405 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_406 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_407 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_408 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_409 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_410 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_411 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_412 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[10]));
 sg13g2_antennanp ANTENNA_413 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[11]));
 sg13g2_antennanp ANTENNA_414 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[12]));
 sg13g2_antennanp ANTENNA_415 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[13]));
 sg13g2_antennanp ANTENNA_416 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[14]));
 sg13g2_antennanp ANTENNA_417 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[15]));
 sg13g2_antennanp ANTENNA_418 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[15]));
 sg13g2_antennanp ANTENNA_419 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[15]));
 sg13g2_antennanp ANTENNA_420 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[16]));
 sg13g2_antennanp ANTENNA_421 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[17]));
 sg13g2_antennanp ANTENNA_422 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[18]));
 sg13g2_antennanp ANTENNA_423 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[19]));
 sg13g2_antennanp ANTENNA_424 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[20]));
 sg13g2_antennanp ANTENNA_425 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[21]));
 sg13g2_antennanp ANTENNA_426 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[22]));
 sg13g2_antennanp ANTENNA_427 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[22]));
 sg13g2_antennanp ANTENNA_428 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[22]));
 sg13g2_antennanp ANTENNA_429 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[23]));
 sg13g2_antennanp ANTENNA_430 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[24]));
 sg13g2_antennanp ANTENNA_431 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[25]));
 sg13g2_antennanp ANTENNA_432 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_433 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[27]));
 sg13g2_antennanp ANTENNA_434 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[28]));
 sg13g2_antennanp ANTENNA_435 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[29]));
 sg13g2_antennanp ANTENNA_436 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[2]));
 sg13g2_antennanp ANTENNA_437 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_438 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[31]));
 sg13g2_antennanp ANTENNA_439 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[3]));
 sg13g2_antennanp ANTENNA_440 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[4]));
 sg13g2_antennanp ANTENNA_441 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[5]));
 sg13g2_antennanp ANTENNA_442 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[6]));
 sg13g2_antennanp ANTENNA_443 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[7]));
 sg13g2_antennanp ANTENNA_444 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[8]));
 sg13g2_antennanp ANTENNA_445 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[9]));
 sg13g2_antennanp ANTENNA_446 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_gnt_i));
 sg13g2_antennanp ANTENNA_447 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[13]));
 sg13g2_antennanp ANTENNA_448 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[13]));
 sg13g2_antennanp ANTENNA_449 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[13]));
 sg13g2_antennanp ANTENNA_450 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[13]));
 sg13g2_antennanp ANTENNA_451 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_452 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_453 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_454 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_455 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_456 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_457 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_458 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_459 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_460 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_461 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_462 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[2]));
 sg13g2_antennanp ANTENNA_463 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_464 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_465 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_466 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_467 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[9]));
 sg13g2_antennanp ANTENNA_468 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[9]));
 sg13g2_antennanp ANTENNA_469 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_470 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_471 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_472 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_473 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_474 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_475 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_476 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_477 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_478 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_479 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_480 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_481 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_482 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_483 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_484 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_485 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[1]));
 sg13g2_antennanp ANTENNA_486 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_busy ));
 sg13g2_antennanp ANTENNA_487 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_488 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_489 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_490 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_491 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/pc_mux_id [1]));
 sg13g2_antennanp ANTENNA_492 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/perf_instr_ret_wb ));
 sg13g2_antennanp ANTENNA_493 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_494 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_495 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_496 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_497 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_498 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_499 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_500 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_501 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_502 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_503 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_504 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_505 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/id_stage_i/_0455_ ));
 sg13g2_antennanp ANTENNA_506 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_507 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_508 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_509 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_510 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_511 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_512 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_148_ ));
 sg13g2_antennanp ANTENNA_513 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_514 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_515 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_516 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_517 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_518 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_519 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_520 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_521 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_522 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_523 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_524 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_525 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_526 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_527 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_528 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_529 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_530 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_531 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_532 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_533 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_534 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_535 (.VDD(VDD),
    .VSS(VSS),
    .A(net1720));
 sg13g2_antennanp ANTENNA_536 (.VDD(VDD),
    .VSS(VSS),
    .A(net1736));
 sg13g2_antennanp ANTENNA_537 (.VDD(VDD),
    .VSS(VSS),
    .A(net1742));
 sg13g2_antennanp ANTENNA_538 (.VDD(VDD),
    .VSS(VSS),
    .A(net1752));
 sg13g2_antennanp ANTENNA_539 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 sg13g2_antennanp ANTENNA_540 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 sg13g2_antennanp ANTENNA_541 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_542 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_543 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_544 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_545 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_546 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_547 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[11]));
 sg13g2_antennanp ANTENNA_548 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_549 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_550 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[13]));
 sg13g2_antennanp ANTENNA_551 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_552 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_553 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[15]));
 sg13g2_antennanp ANTENNA_554 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[16]));
 sg13g2_antennanp ANTENNA_555 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[16]));
 sg13g2_antennanp ANTENNA_556 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[17]));
 sg13g2_antennanp ANTENNA_557 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[18]));
 sg13g2_antennanp ANTENNA_558 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[19]));
 sg13g2_antennanp ANTENNA_559 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[19]));
 sg13g2_antennanp ANTENNA_560 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[20]));
 sg13g2_antennanp ANTENNA_561 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[21]));
 sg13g2_antennanp ANTENNA_562 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[23]));
 sg13g2_antennanp ANTENNA_563 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_564 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_565 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[25]));
 sg13g2_antennanp ANTENNA_566 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_567 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_568 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[27]));
 sg13g2_antennanp ANTENNA_569 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[28]));
 sg13g2_antennanp ANTENNA_570 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[29]));
 sg13g2_antennanp ANTENNA_571 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_572 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_573 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[31]));
 sg13g2_antennanp ANTENNA_574 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[9]));
 sg13g2_antennanp ANTENNA_575 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_576 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_577 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_578 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_579 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_580 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_581 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_582 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_583 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_584 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_585 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_586 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_587 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_588 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_589 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_590 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_591 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_592 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_593 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_594 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_595 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_596 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_597 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_598 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_599 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_600 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_601 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_602 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_603 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_604 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_605 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_606 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_607 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_608 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_609 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_610 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_611 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_612 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_613 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[17]));
 sg13g2_antennanp ANTENNA_614 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_615 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_616 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_617 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_618 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_619 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_620 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_621 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_622 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_623 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_624 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_625 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_626 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_627 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_628 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_629 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_630 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_631 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_632 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_633 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_634 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_635 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_636 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_637 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_638 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_639 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_640 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_641 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_642 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_643 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_644 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_645 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_646 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_647 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_648 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_649 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_650 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_651 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_652 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_653 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_654 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_655 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_656 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_657 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_658 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_659 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[10]));
 sg13g2_antennanp ANTENNA_660 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[11]));
 sg13g2_antennanp ANTENNA_661 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[12]));
 sg13g2_antennanp ANTENNA_662 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[13]));
 sg13g2_antennanp ANTENNA_663 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[14]));
 sg13g2_antennanp ANTENNA_664 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[15]));
 sg13g2_antennanp ANTENNA_665 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[16]));
 sg13g2_antennanp ANTENNA_666 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[17]));
 sg13g2_antennanp ANTENNA_667 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[18]));
 sg13g2_antennanp ANTENNA_668 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[19]));
 sg13g2_antennanp ANTENNA_669 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[20]));
 sg13g2_antennanp ANTENNA_670 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[21]));
 sg13g2_antennanp ANTENNA_671 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[22]));
 sg13g2_antennanp ANTENNA_672 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[23]));
 sg13g2_antennanp ANTENNA_673 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[24]));
 sg13g2_antennanp ANTENNA_674 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[25]));
 sg13g2_antennanp ANTENNA_675 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_676 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_677 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_678 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[27]));
 sg13g2_antennanp ANTENNA_679 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[28]));
 sg13g2_antennanp ANTENNA_680 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[29]));
 sg13g2_antennanp ANTENNA_681 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[2]));
 sg13g2_antennanp ANTENNA_682 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[2]));
 sg13g2_antennanp ANTENNA_683 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[2]));
 sg13g2_antennanp ANTENNA_684 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_685 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_686 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_687 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[31]));
 sg13g2_antennanp ANTENNA_688 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[3]));
 sg13g2_antennanp ANTENNA_689 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[4]));
 sg13g2_antennanp ANTENNA_690 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[5]));
 sg13g2_antennanp ANTENNA_691 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[6]));
 sg13g2_antennanp ANTENNA_692 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[7]));
 sg13g2_antennanp ANTENNA_693 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[8]));
 sg13g2_antennanp ANTENNA_694 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[9]));
 sg13g2_antennanp ANTENNA_695 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_gnt_i));
 sg13g2_antennanp ANTENNA_696 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_697 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_698 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_699 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_700 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_701 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_702 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_703 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_704 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_705 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_706 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_707 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[2]));
 sg13g2_antennanp ANTENNA_708 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_709 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_710 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_711 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_712 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_713 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_714 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_715 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_716 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_717 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_busy ));
 sg13g2_antennanp ANTENNA_718 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_719 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_720 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_721 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_722 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/pc_mux_id [1]));
 sg13g2_antennanp ANTENNA_723 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/perf_instr_ret_wb ));
 sg13g2_antennanp ANTENNA_724 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_725 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_726 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_727 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_728 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_729 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_730 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_731 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_732 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_733 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_734 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_735 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_736 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/id_stage_i/_0455_ ));
 sg13g2_antennanp ANTENNA_737 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_738 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_739 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_740 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_741 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_742 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_743 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_744 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_745 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_746 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_747 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_748 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_749 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_750 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_751 (.VDD(VDD),
    .VSS(VSS),
    .A(net1720));
 sg13g2_antennanp ANTENNA_752 (.VDD(VDD),
    .VSS(VSS),
    .A(net1742));
 sg13g2_antennanp ANTENNA_753 (.VDD(VDD),
    .VSS(VSS),
    .A(net1752));
 sg13g2_antennanp ANTENNA_754 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 sg13g2_antennanp ANTENNA_755 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 sg13g2_antennanp ANTENNA_756 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_757 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_758 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_759 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_760 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_761 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_762 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[10]));
 sg13g2_antennanp ANTENNA_763 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[11]));
 sg13g2_antennanp ANTENNA_764 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_765 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[12]));
 sg13g2_antennanp ANTENNA_766 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[13]));
 sg13g2_antennanp ANTENNA_767 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_768 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[14]));
 sg13g2_antennanp ANTENNA_769 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[15]));
 sg13g2_antennanp ANTENNA_770 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[16]));
 sg13g2_antennanp ANTENNA_771 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[17]));
 sg13g2_antennanp ANTENNA_772 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[18]));
 sg13g2_antennanp ANTENNA_773 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[19]));
 sg13g2_antennanp ANTENNA_774 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[19]));
 sg13g2_antennanp ANTENNA_775 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[20]));
 sg13g2_antennanp ANTENNA_776 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[21]));
 sg13g2_antennanp ANTENNA_777 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[23]));
 sg13g2_antennanp ANTENNA_778 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_779 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[24]));
 sg13g2_antennanp ANTENNA_780 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[25]));
 sg13g2_antennanp ANTENNA_781 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_782 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[26]));
 sg13g2_antennanp ANTENNA_783 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[27]));
 sg13g2_antennanp ANTENNA_784 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[28]));
 sg13g2_antennanp ANTENNA_785 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[29]));
 sg13g2_antennanp ANTENNA_786 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_787 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[30]));
 sg13g2_antennanp ANTENNA_788 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[31]));
 sg13g2_antennanp ANTENNA_789 (.VDD(VDD),
    .VSS(VSS),
    .A(boot_addr_i[9]));
 sg13g2_antennanp ANTENNA_790 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_791 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_792 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_793 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_794 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_795 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_796 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[11]));
 sg13g2_antennanp ANTENNA_797 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_798 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_799 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_800 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_801 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_802 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[12]));
 sg13g2_antennanp ANTENNA_803 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_804 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_805 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_806 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_807 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_808 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_809 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[13]));
 sg13g2_antennanp ANTENNA_810 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_811 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_812 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_813 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_814 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_815 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_816 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[14]));
 sg13g2_antennanp ANTENNA_817 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_818 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_819 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_820 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_821 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_822 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[16]));
 sg13g2_antennanp ANTENNA_823 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_824 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_825 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_826 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_827 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_828 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_829 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[19]));
 sg13g2_antennanp ANTENNA_830 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_831 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_832 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_833 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_834 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_835 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_836 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[20]));
 sg13g2_antennanp ANTENNA_837 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_838 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_839 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_840 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_841 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_842 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_843 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[21]));
 sg13g2_antennanp ANTENNA_844 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_845 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_846 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_847 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_848 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_849 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[22]));
 sg13g2_antennanp ANTENNA_850 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_851 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_852 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_853 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_854 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[25]));
 sg13g2_antennanp ANTENNA_855 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_856 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_857 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_858 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_859 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[27]));
 sg13g2_antennanp ANTENNA_860 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_861 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_862 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_863 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_864 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_865 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_866 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_867 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_868 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[28]));
 sg13g2_antennanp ANTENNA_869 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_870 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_871 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_872 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_873 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[30]));
 sg13g2_antennanp ANTENNA_874 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_875 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_876 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_877 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_878 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_879 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_880 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[8]));
 sg13g2_antennanp ANTENNA_881 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_882 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_883 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_884 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_885 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_886 (.VDD(VDD),
    .VSS(VSS),
    .A(data_rdata_i[9]));
 sg13g2_antennanp ANTENNA_887 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_888 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_889 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_890 (.VDD(VDD),
    .VSS(VSS),
    .A(debug_req_i));
 sg13g2_antennanp ANTENNA_891 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[10]));
 sg13g2_antennanp ANTENNA_892 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[11]));
 sg13g2_antennanp ANTENNA_893 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[12]));
 sg13g2_antennanp ANTENNA_894 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[13]));
 sg13g2_antennanp ANTENNA_895 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[14]));
 sg13g2_antennanp ANTENNA_896 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[15]));
 sg13g2_antennanp ANTENNA_897 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[16]));
 sg13g2_antennanp ANTENNA_898 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[17]));
 sg13g2_antennanp ANTENNA_899 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[18]));
 sg13g2_antennanp ANTENNA_900 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[19]));
 sg13g2_antennanp ANTENNA_901 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[20]));
 sg13g2_antennanp ANTENNA_902 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[21]));
 sg13g2_antennanp ANTENNA_903 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[22]));
 sg13g2_antennanp ANTENNA_904 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[23]));
 sg13g2_antennanp ANTENNA_905 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[24]));
 sg13g2_antennanp ANTENNA_906 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[25]));
 sg13g2_antennanp ANTENNA_907 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_908 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_909 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[26]));
 sg13g2_antennanp ANTENNA_910 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[27]));
 sg13g2_antennanp ANTENNA_911 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[28]));
 sg13g2_antennanp ANTENNA_912 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[29]));
 sg13g2_antennanp ANTENNA_913 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[2]));
 sg13g2_antennanp ANTENNA_914 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_915 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_916 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[30]));
 sg13g2_antennanp ANTENNA_917 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[31]));
 sg13g2_antennanp ANTENNA_918 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[3]));
 sg13g2_antennanp ANTENNA_919 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[4]));
 sg13g2_antennanp ANTENNA_920 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[5]));
 sg13g2_antennanp ANTENNA_921 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[5]));
 sg13g2_antennanp ANTENNA_922 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[5]));
 sg13g2_antennanp ANTENNA_923 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[6]));
 sg13g2_antennanp ANTENNA_924 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[7]));
 sg13g2_antennanp ANTENNA_925 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[8]));
 sg13g2_antennanp ANTENNA_926 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_addr_o[9]));
 sg13g2_antennanp ANTENNA_927 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_gnt_i));
 sg13g2_antennanp ANTENNA_928 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_929 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_930 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_931 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[1]));
 sg13g2_antennanp ANTENNA_932 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_933 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_934 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_935 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_936 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[23]));
 sg13g2_antennanp ANTENNA_937 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_938 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[25]));
 sg13g2_antennanp ANTENNA_939 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[2]));
 sg13g2_antennanp ANTENNA_940 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_941 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[30]));
 sg13g2_antennanp ANTENNA_942 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_943 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rdata_i[5]));
 sg13g2_antennanp ANTENNA_944 (.VDD(VDD),
    .VSS(VSS),
    .A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_945 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_946 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_947 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_948 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[11]));
 sg13g2_antennanp ANTENNA_949 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_950 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_951 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_952 (.VDD(VDD),
    .VSS(VSS),
    .A(irqs_i[15]));
 sg13g2_antennanp ANTENNA_953 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_busy ));
 sg13g2_antennanp ANTENNA_954 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_955 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_956 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_957 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/instr_req_gated ));
 sg13g2_antennanp ANTENNA_958 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/pc_mux_id [1]));
 sg13g2_antennanp ANTENNA_959 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/perf_instr_ret_wb ));
 sg13g2_antennanp ANTENNA_960 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_961 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/cs_registers_i/minstret_counter_i/_0077_ ));
 sg13g2_antennanp ANTENNA_962 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_963 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_964 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_965 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_966 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_967 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_968 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_969 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_970 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_971 (.VDD(VDD),
    .VSS(VSS),
    .A(net698));
 sg13g2_antennanp ANTENNA_972 (.VDD(VDD),
    .VSS(VSS),
    .A(\i_ibex/if_stage_i/prefetch_buffer_i/fifo_i/_225_ ));
 sg13g2_antennanp ANTENNA_973 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_974 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_975 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_976 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_977 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_978 (.VDD(VDD),
    .VSS(VSS),
    .A(net1484));
 sg13g2_antennanp ANTENNA_979 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_980 (.VDD(VDD),
    .VSS(VSS),
    .A(net1500));
 sg13g2_antennanp ANTENNA_981 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_982 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_983 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_984 (.VDD(VDD),
    .VSS(VSS),
    .A(net1502));
 sg13g2_antennanp ANTENNA_985 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_986 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_987 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_988 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_989 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_990 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_991 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_992 (.VDD(VDD),
    .VSS(VSS),
    .A(net1581));
 sg13g2_antennanp ANTENNA_993 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_994 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_995 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_996 (.VDD(VDD),
    .VSS(VSS),
    .A(net1613));
 sg13g2_antennanp ANTENNA_997 (.VDD(VDD),
    .VSS(VSS),
    .A(net1720));
 sg13g2_antennanp ANTENNA_998 (.VDD(VDD),
    .VSS(VSS),
    .A(net1742));
 sg13g2_antennanp ANTENNA_999 (.VDD(VDD),
    .VSS(VSS),
    .A(net1752));
 sg13g2_antennanp ANTENNA_1000 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 sg13g2_antennanp ANTENNA_1001 (.VDD(VDD),
    .VSS(VSS),
    .A(net1767));
 assign data_addr_o[1] = data_addr_o[0];
 assign instr_addr_o[1] = instr_addr_o[0];
endmodule
