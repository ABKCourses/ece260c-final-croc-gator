module cve2_register_file_ff (clk_i,
    rst_ni,
    test_en_i,
    we_a_i,
    raddr_a_i,
    raddr_b_i,
    rdata_a_o,
    rdata_b_o,
    waddr_a_i,
    wdata_a_i);
 input clk_i;
 input rst_ni;
 input test_en_i;
 input we_a_i;
 input [4:0] raddr_a_i;
 input [4:0] raddr_b_i;
 output [31:0] rdata_a_o;
 output [31:0] rdata_b_o;
 input [4:0] waddr_a_i;
 input [31:0] wdata_a_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire clknet_leaf_33_clk_i;
 wire _0993_;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_27_clk_i;
 wire _1000_;
 wire clknet_leaf_26_clk_i;
 wire _1002_;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_22_clk_i;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_20_clk_i;
 wire _1013_;
 wire _1014_;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_18_clk_i;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire clknet_leaf_17_clk_i;
 wire _1021_;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_13_clk_i;
 wire _1026_;
 wire _1027_;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_7_clk_i;
 wire _1034_;
 wire clknet_leaf_6_clk_i;
 wire _1036_;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_4_clk_i;
 wire _1039_;
 wire clknet_leaf_3_clk_i;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire clknet_leaf_2_clk_i;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_0_clk_i;
 wire _1051_;
 wire _1052_;
 wire net315;
 wire _1054_;
 wire net314;
 wire net313;
 wire _1057_;
 wire net312;
 wire _1059_;
 wire net311;
 wire _1061_;
 wire net310;
 wire net309;
 wire _1064_;
 wire net308;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire net307;
 wire _1073_;
 wire net306;
 wire _1075_;
 wire net305;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire net304;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire net303;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire net302;
 wire net301;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire net300;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire net299;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire net298;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire net297;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire net296;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire net295;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire net294;
 wire _1233_;
 wire _1234_;
 wire net293;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire net292;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire net291;
 wire _1261_;
 wire _1262_;
 wire net290;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire net289;
 wire _1281_;
 wire _1282_;
 wire net288;
 wire _1284_;
 wire _1285_;
 wire net287;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire net286;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire net285;
 wire net284;
 wire _1298_;
 wire _1299_;
 wire net283;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire net282;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire net281;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire net280;
 wire _1337_;
 wire net279;
 wire _1339_;
 wire _1340_;
 wire net278;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire net277;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire net276;
 wire _1352_;
 wire net275;
 wire _1354_;
 wire _1355_;
 wire net274;
 wire net273;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire net272;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire net271;
 wire _1370_;
 wire net270;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire net269;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire net268;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire net267;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire net266;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire net265;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire net264;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire net263;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire net262;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire net261;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire net260;
 wire _1527_;
 wire _1528_;
 wire net259;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire net258;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire net257;
 wire _1555_;
 wire _1556_;
 wire net256;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire net255;
 wire _1575_;
 wire _1576_;
 wire net254;
 wire _1578_;
 wire _1579_;
 wire net253;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire net252;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire net251;
 wire net250;
 wire _1592_;
 wire _1593_;
 wire net249;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire net248;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire net247;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire net246;
 wire _1631_;
 wire net245;
 wire _1633_;
 wire _1634_;
 wire net244;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire net243;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire net242;
 wire _1646_;
 wire net241;
 wire _1648_;
 wire _1649_;
 wire net240;
 wire net239;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire net238;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire net237;
 wire _1664_;
 wire net236;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire net235;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire net234;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire net233;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire net232;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire net231;
 wire net230;
 wire net229;
 wire net228;
 wire net227;
 wire net226;
 wire net225;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire net224;
 wire net223;
 wire net222;
 wire net221;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire net220;
 wire net219;
 wire net218;
 wire net217;
 wire net216;
 wire net215;
 wire _1979_;
 wire net214;
 wire net213;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire net212;
 wire _1986_;
 wire net211;
 wire net210;
 wire _1989_;
 wire net209;
 wire net208;
 wire _1992_;
 wire _1993_;
 wire net207;
 wire net206;
 wire net205;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire net204;
 wire net203;
 wire _2002_;
 wire net202;
 wire net201;
 wire _2005_;
 wire _2006_;
 wire net200;
 wire net199;
 wire _2009_;
 wire _2010_;
 wire net198;
 wire net197;
 wire _2013_;
 wire _2014_;
 wire net196;
 wire net195;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire net194;
 wire _2021_;
 wire net193;
 wire _2023_;
 wire net192;
 wire _2025_;
 wire net191;
 wire net190;
 wire _2028_;
 wire net189;
 wire _2030_;
 wire net188;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire net187;
 wire net186;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire net185;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire net184;
 wire _2052_;
 wire net183;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire net182;
 wire net181;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire net180;
 wire _2120_;
 wire net179;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire net178;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire net177;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire net176;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire net175;
 wire _2172_;
 wire net174;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire net173;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire net172;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire net171;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire net170;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire net169;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire net168;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire net167;
 wire net166;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire net165;
 wire _2265_;
 wire _2266_;
 wire net164;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire net163;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire net162;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire net161;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire net160;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire net159;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire net158;
 wire net157;
 wire net156;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire net155;
 wire _2319_;
 wire _2320_;
 wire net154;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire net153;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire net152;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire net151;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire net150;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire net149;
 wire _2357_;
 wire net148;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire net147;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire net146;
 wire _2424_;
 wire net145;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire net144;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire net143;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire net142;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire net141;
 wire _2476_;
 wire net140;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire net139;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire net138;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire net137;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire net136;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire net135;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire net134;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire net133;
 wire net132;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire net131;
 wire _2569_;
 wire _2570_;
 wire net130;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire net129;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire net128;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire net127;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire net126;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire net125;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire net124;
 wire net123;
 wire net122;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire net121;
 wire _2623_;
 wire _2624_;
 wire net120;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire net119;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire net118;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire net117;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire net116;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire net115;
 wire _2661_;
 wire net114;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire net113;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire net112;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire net111;
 wire net110;
 wire net109;
 wire net108;
 wire net107;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire _2963_;
 wire net100;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire _3016_;
 wire net52;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire _3028_;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire _3037_;
 wire _3038_;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire _3045_;
 wire net30;
 wire net29;
 wire net28;
 wire _3049_;
 wire net27;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire _3058_;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire _3063_;
 wire net18;
 wire _3065_;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire _3070_;
 wire net13;
 wire net12;
 wire net11;
 wire _3074_;
 wire net10;
 wire net9;
 wire net8;
 wire _3078_;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire _3083_;
 wire net3;
 wire net2;
 wire net1;
 wire _3087_;
 wire clknet_leaf_122_clk_i;
 wire clknet_leaf_121_clk_i;
 wire clknet_leaf_120_clk_i;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire clknet_leaf_119_clk_i;
 wire clknet_leaf_118_clk_i;
 wire clknet_leaf_117_clk_i;
 wire clknet_leaf_116_clk_i;
 wire clknet_leaf_115_clk_i;
 wire _3099_;
 wire clknet_leaf_114_clk_i;
 wire clknet_leaf_113_clk_i;
 wire clknet_leaf_112_clk_i;
 wire clknet_leaf_111_clk_i;
 wire _3104_;
 wire _3105_;
 wire clknet_leaf_110_clk_i;
 wire clknet_leaf_109_clk_i;
 wire clknet_leaf_108_clk_i;
 wire clknet_leaf_107_clk_i;
 wire clknet_leaf_106_clk_i;
 wire clknet_leaf_105_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_90_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_85_clk_i;
 wire clknet_leaf_84_clk_i;
 wire _3133_;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_82_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_80_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_76_clk_i;
 wire _3142_;
 wire _3143_;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_72_clk_i;
 wire _3148_;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_68_clk_i;
 wire _3153_;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_65_clk_i;
 wire _3157_;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_62_clk_i;
 wire _3161_;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_58_clk_i;
 wire _3166_;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_55_clk_i;
 wire clknet_leaf_54_clk_i;
 wire _3171_;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_50_clk_i;
 wire _3176_;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_46_clk_i;
 wire _3181_;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_43_clk_i;
 wire _3185_;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_40_clk_i;
 wire _3189_;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_37_clk_i;
 wire _3193_;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_34_clk_i;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire clknet_leaf_123_clk_i;
 wire VDD;
 wire VSS;
 wire clknet_leaf_124_clk_i;
 wire clknet_leaf_125_clk_i;
 wire clknet_leaf_126_clk_i;
 wire clknet_leaf_127_clk_i;
 wire clknet_leaf_128_clk_i;
 wire clknet_leaf_129_clk_i;
 wire clknet_leaf_130_clk_i;
 wire clknet_0_clk_i;
 wire clknet_4_0_0_clk_i;
 wire clknet_4_1_0_clk_i;
 wire clknet_4_2_0_clk_i;
 wire clknet_4_3_0_clk_i;
 wire clknet_4_4_0_clk_i;
 wire clknet_4_5_0_clk_i;
 wire clknet_4_6_0_clk_i;
 wire clknet_4_7_0_clk_i;
 wire clknet_4_8_0_clk_i;
 wire clknet_4_9_0_clk_i;
 wire clknet_4_10_0_clk_i;
 wire clknet_4_11_0_clk_i;
 wire clknet_4_12_0_clk_i;
 wire clknet_4_13_0_clk_i;
 wire clknet_4_14_0_clk_i;
 wire clknet_4_15_0_clk_i;
 wire clknet_5_0__leaf_clk_i;
 wire clknet_5_1__leaf_clk_i;
 wire clknet_5_2__leaf_clk_i;
 wire clknet_5_3__leaf_clk_i;
 wire clknet_5_4__leaf_clk_i;
 wire clknet_5_5__leaf_clk_i;
 wire clknet_5_6__leaf_clk_i;
 wire clknet_5_7__leaf_clk_i;
 wire clknet_5_8__leaf_clk_i;
 wire clknet_5_9__leaf_clk_i;
 wire clknet_5_10__leaf_clk_i;
 wire clknet_5_11__leaf_clk_i;
 wire clknet_5_12__leaf_clk_i;
 wire clknet_5_13__leaf_clk_i;
 wire clknet_5_14__leaf_clk_i;
 wire clknet_5_15__leaf_clk_i;
 wire clknet_5_16__leaf_clk_i;
 wire clknet_5_17__leaf_clk_i;
 wire clknet_5_18__leaf_clk_i;
 wire clknet_5_19__leaf_clk_i;
 wire clknet_5_20__leaf_clk_i;
 wire clknet_5_21__leaf_clk_i;
 wire clknet_5_22__leaf_clk_i;
 wire clknet_5_23__leaf_clk_i;
 wire clknet_5_24__leaf_clk_i;
 wire clknet_5_25__leaf_clk_i;
 wire clknet_5_26__leaf_clk_i;
 wire clknet_5_27__leaf_clk_i;
 wire clknet_5_28__leaf_clk_i;
 wire clknet_5_29__leaf_clk_i;
 wire clknet_5_30__leaf_clk_i;
 wire clknet_5_31__leaf_clk_i;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire [1023:0] rf_reg;

 sg13g2_mux2_1 _4190_ (.A0(rf_reg[477]),
    .A1(net335),
    .S(net1),
    .X(_0416_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4191_ (.A0(rf_reg[478]),
    .A1(net319),
    .S(net2),
    .X(_0417_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4192_ (.A0(rf_reg[479]),
    .A1(net323),
    .S(net2),
    .X(_0418_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4193_ (.A0(net332),
    .A1(rf_reg[47]),
    .S(net25),
    .X(_0419_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4194_ (.A(_2949_),
    .B(_3037_),
    .Y(_3087_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_122_clk_i (.X(clknet_leaf_122_clk_i),
    .A(clknet_5_5__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4196_ (.A0(rf_reg[480]),
    .A1(net328),
    .S(net154),
    .X(_0420_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4197_ (.A0(rf_reg[481]),
    .A1(net329),
    .S(net154),
    .X(_0421_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4198_ (.A0(rf_reg[482]),
    .A1(net346),
    .S(net151),
    .X(_0422_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4199_ (.A0(rf_reg[483]),
    .A1(net331),
    .S(net153),
    .X(_0423_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4200_ (.A0(rf_reg[484]),
    .A1(net337),
    .S(net151),
    .X(_0424_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4201_ (.A0(rf_reg[485]),
    .A1(net342),
    .S(net153),
    .X(_0425_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4202_ (.A0(rf_reg[486]),
    .A1(net326),
    .S(net152),
    .X(_0426_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4203_ (.A0(rf_reg[487]),
    .A1(net340),
    .S(net153),
    .X(_0427_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4204_ (.A0(rf_reg[488]),
    .A1(net341),
    .S(net151),
    .X(_0428_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4205_ (.A0(rf_reg[489]),
    .A1(net347),
    .S(net151),
    .X(_0429_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4206_ (.A0(net320),
    .A1(rf_reg[48]),
    .S(net25),
    .X(_0430_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_121_clk_i (.X(clknet_leaf_121_clk_i),
    .A(clknet_5_5__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4208_ (.A0(rf_reg[490]),
    .A1(net327),
    .S(net152),
    .X(_0431_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4209_ (.A0(rf_reg[491]),
    .A1(net317),
    .S(net154),
    .X(_0432_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4210_ (.A0(rf_reg[492]),
    .A1(net322),
    .S(net152),
    .X(_0433_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4211_ (.A0(rf_reg[493]),
    .A1(net345),
    .S(net153),
    .X(_0434_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4212_ (.A0(rf_reg[494]),
    .A1(net321),
    .S(net152),
    .X(_0435_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4213_ (.A0(rf_reg[495]),
    .A1(net332),
    .S(net154),
    .X(_0436_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4214_ (.A0(rf_reg[496]),
    .A1(net320),
    .S(net154),
    .X(_0437_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4215_ (.A0(rf_reg[497]),
    .A1(net330),
    .S(net151),
    .X(_0438_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4216_ (.A0(rf_reg[498]),
    .A1(net318),
    .S(net154),
    .X(_0439_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4217_ (.A0(rf_reg[499]),
    .A1(net325),
    .S(net154),
    .X(_0440_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4218_ (.A0(net330),
    .A1(rf_reg[49]),
    .S(net22),
    .X(_0441_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_120_clk_i (.X(clknet_leaf_120_clk_i),
    .A(clknet_5_5__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4220_ (.A0(rf_reg[500]),
    .A1(net344),
    .S(net153),
    .X(_0442_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4221_ (.A0(rf_reg[501]),
    .A1(net334),
    .S(net152),
    .X(_0443_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4222_ (.A0(rf_reg[502]),
    .A1(net338),
    .S(net151),
    .X(_0444_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4223_ (.A0(rf_reg[503]),
    .A1(net324),
    .S(net155),
    .X(_0445_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4224_ (.A0(rf_reg[504]),
    .A1(net336),
    .S(net153),
    .X(_0446_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4225_ (.A0(rf_reg[505]),
    .A1(net333),
    .S(net155),
    .X(_0447_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4226_ (.A0(rf_reg[506]),
    .A1(net343),
    .S(net151),
    .X(_0448_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4227_ (.A0(rf_reg[507]),
    .A1(net316),
    .S(net153),
    .X(_0449_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4228_ (.A0(rf_reg[508]),
    .A1(net339),
    .S(net153),
    .X(_0450_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4229_ (.A0(rf_reg[509]),
    .A1(net335),
    .S(net151),
    .X(_0451_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4230_ (.A0(net318),
    .A1(rf_reg[50]),
    .S(net24),
    .X(_0452_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4231_ (.A0(rf_reg[510]),
    .A1(net319),
    .S(net152),
    .X(_0453_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4232_ (.A0(rf_reg[511]),
    .A1(net323),
    .S(net152),
    .X(_0454_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _4233_ (.Y(_3091_),
    .A(waddr_a_i[4]),
    .B(we_a_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 _4234_ (.A(_3091_),
    .B_N(_3051_),
    .Y(_3092_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _4235_ (.Y(_3093_),
    .B(_3092_),
    .A_N(_3016_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_119_clk_i (.X(clknet_leaf_119_clk_i),
    .A(clknet_5_4__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_118_clk_i (.X(clknet_leaf_118_clk_i),
    .A(clknet_5_6__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4238_ (.A0(net328),
    .A1(rf_reg[512]),
    .S(net148),
    .X(_0455_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4239_ (.A0(net329),
    .A1(rf_reg[513]),
    .S(net148),
    .X(_0456_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4240_ (.A0(net346),
    .A1(rf_reg[514]),
    .S(net146),
    .X(_0457_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4241_ (.A0(net331),
    .A1(rf_reg[515]),
    .S(net149),
    .X(_0458_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4242_ (.A0(net337),
    .A1(rf_reg[516]),
    .S(net147),
    .X(_0459_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4243_ (.A0(net342),
    .A1(rf_reg[517]),
    .S(net149),
    .X(_0460_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4244_ (.A0(net326),
    .A1(rf_reg[518]),
    .S(net146),
    .X(_0461_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4245_ (.A0(net340),
    .A1(rf_reg[519]),
    .S(net148),
    .X(_0462_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4246_ (.A0(net325),
    .A1(rf_reg[51]),
    .S(net24),
    .X(_0463_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4247_ (.A0(net341),
    .A1(rf_reg[520]),
    .S(net146),
    .X(_0464_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4248_ (.A0(net347),
    .A1(rf_reg[521]),
    .S(net146),
    .X(_0465_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_117_clk_i (.X(clknet_leaf_117_clk_i),
    .A(clknet_5_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4250_ (.A0(net327),
    .A1(rf_reg[522]),
    .S(net150),
    .X(_0466_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4251_ (.A0(net317),
    .A1(rf_reg[523]),
    .S(net148),
    .X(_0467_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4252_ (.A0(net322),
    .A1(rf_reg[524]),
    .S(net147),
    .X(_0468_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4253_ (.A0(net345),
    .A1(rf_reg[525]),
    .S(net149),
    .X(_0469_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4254_ (.A0(net321),
    .A1(rf_reg[526]),
    .S(net147),
    .X(_0470_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4255_ (.A0(net332),
    .A1(rf_reg[527]),
    .S(net147),
    .X(_0471_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4256_ (.A0(net320),
    .A1(rf_reg[528]),
    .S(net148),
    .X(_0472_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4257_ (.A0(net330),
    .A1(rf_reg[529]),
    .S(net146),
    .X(_0473_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_116_clk_i (.X(clknet_leaf_116_clk_i),
    .A(clknet_5_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4259_ (.A0(net344),
    .A1(rf_reg[52]),
    .S(net23),
    .X(_0474_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4260_ (.A0(net318),
    .A1(rf_reg[530]),
    .S(net148),
    .X(_0475_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4261_ (.A0(net325),
    .A1(rf_reg[531]),
    .S(net148),
    .X(_0476_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_115_clk_i (.X(clknet_leaf_115_clk_i),
    .A(clknet_5_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4263_ (.A0(net344),
    .A1(rf_reg[532]),
    .S(net149),
    .X(_0477_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4264_ (.A0(net334),
    .A1(rf_reg[533]),
    .S(net146),
    .X(_0478_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4265_ (.A0(net338),
    .A1(rf_reg[534]),
    .S(net146),
    .X(_0479_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4266_ (.A0(net324),
    .A1(rf_reg[535]),
    .S(net149),
    .X(_0480_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4267_ (.A0(net336),
    .A1(rf_reg[536]),
    .S(net149),
    .X(_0481_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4268_ (.A0(net333),
    .A1(rf_reg[537]),
    .S(net150),
    .X(_0482_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4269_ (.A0(net343),
    .A1(rf_reg[538]),
    .S(net147),
    .X(_0483_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4270_ (.A0(net316),
    .A1(rf_reg[539]),
    .S(net148),
    .X(_0484_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4271_ (.A0(net334),
    .A1(rf_reg[53]),
    .S(net21),
    .X(_0485_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4272_ (.A0(net339),
    .A1(rf_reg[540]),
    .S(net149),
    .X(_0486_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4273_ (.A0(net335),
    .A1(rf_reg[541]),
    .S(net146),
    .X(_0487_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4274_ (.A0(net319),
    .A1(rf_reg[542]),
    .S(net147),
    .X(_0488_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4275_ (.A0(net323),
    .A1(rf_reg[543]),
    .S(net147),
    .X(_0489_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _4276_ (.Y(_3099_),
    .B(_3092_),
    .A_N(_2963_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_114_clk_i (.X(clknet_leaf_114_clk_i),
    .A(clknet_5_18__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_113_clk_i (.X(clknet_leaf_113_clk_i),
    .A(clknet_5_18__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4279_ (.A0(net328),
    .A1(rf_reg[544]),
    .S(net143),
    .X(_0490_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4280_ (.A0(net329),
    .A1(rf_reg[545]),
    .S(net143),
    .X(_0491_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4281_ (.A0(net346),
    .A1(rf_reg[546]),
    .S(net141),
    .X(_0492_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4282_ (.A0(net331),
    .A1(rf_reg[547]),
    .S(net144),
    .X(_0493_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4283_ (.A0(net337),
    .A1(rf_reg[548]),
    .S(net142),
    .X(_0494_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4284_ (.A0(net342),
    .A1(rf_reg[549]),
    .S(net144),
    .X(_0495_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4285_ (.A0(net338),
    .A1(rf_reg[54]),
    .S(net21),
    .X(_0496_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4286_ (.A0(net326),
    .A1(rf_reg[550]),
    .S(net142),
    .X(_0497_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4287_ (.A0(net340),
    .A1(rf_reg[551]),
    .S(net144),
    .X(_0498_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4288_ (.A0(net341),
    .A1(rf_reg[552]),
    .S(net141),
    .X(_0499_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4289_ (.A0(net347),
    .A1(rf_reg[553]),
    .S(net141),
    .X(_0500_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_112_clk_i (.X(clknet_leaf_112_clk_i),
    .A(clknet_5_18__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4291_ (.A0(net327),
    .A1(rf_reg[554]),
    .S(net145),
    .X(_0501_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4292_ (.A0(net317),
    .A1(rf_reg[555]),
    .S(net143),
    .X(_0502_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4293_ (.A0(net322),
    .A1(rf_reg[556]),
    .S(net142),
    .X(_0503_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4294_ (.A0(net345),
    .A1(rf_reg[557]),
    .S(net144),
    .X(_0504_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4295_ (.A0(net321),
    .A1(rf_reg[558]),
    .S(net142),
    .X(_0505_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4296_ (.A0(net332),
    .A1(rf_reg[559]),
    .S(net142),
    .X(_0506_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4297_ (.A0(net324),
    .A1(rf_reg[55]),
    .S(net23),
    .X(_0507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4298_ (.A0(net320),
    .A1(rf_reg[560]),
    .S(net143),
    .X(_0508_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4299_ (.A0(net330),
    .A1(rf_reg[561]),
    .S(net141),
    .X(_0509_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4300_ (.A0(net318),
    .A1(rf_reg[562]),
    .S(net143),
    .X(_0510_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4301_ (.A0(net325),
    .A1(rf_reg[563]),
    .S(net143),
    .X(_0511_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_111_clk_i (.X(clknet_leaf_111_clk_i),
    .A(clknet_5_19__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4303_ (.A0(net344),
    .A1(rf_reg[564]),
    .S(net144),
    .X(_0512_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4304_ (.A0(net334),
    .A1(rf_reg[565]),
    .S(net141),
    .X(_0513_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4305_ (.A0(net338),
    .A1(rf_reg[566]),
    .S(net141),
    .X(_0514_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4306_ (.A0(net324),
    .A1(rf_reg[567]),
    .S(net144),
    .X(_0515_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4307_ (.A0(net336),
    .A1(rf_reg[568]),
    .S(net143),
    .X(_0516_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4308_ (.A0(net333),
    .A1(rf_reg[569]),
    .S(net145),
    .X(_0517_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4309_ (.A0(net336),
    .A1(rf_reg[56]),
    .S(net23),
    .X(_0518_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4310_ (.A0(net343),
    .A1(rf_reg[570]),
    .S(net142),
    .X(_0519_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4311_ (.A0(net316),
    .A1(rf_reg[571]),
    .S(net143),
    .X(_0520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4312_ (.A0(net339),
    .A1(rf_reg[572]),
    .S(net144),
    .X(_0521_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4313_ (.A0(net335),
    .A1(rf_reg[573]),
    .S(net141),
    .X(_0522_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4314_ (.A0(net319),
    .A1(rf_reg[574]),
    .S(net142),
    .X(_0523_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4315_ (.A0(net323),
    .A1(rf_reg[575]),
    .S(net141),
    .X(_0524_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 _4316_ (.Y(_3104_),
    .B(_2966_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(_3091_));
 sg13g2_nor2_1 _4317_ (.A(_3016_),
    .B(_3104_),
    .Y(_3105_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_110_clk_i (.X(clknet_leaf_110_clk_i),
    .A(clknet_5_17__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4319_ (.A0(rf_reg[576]),
    .A1(net328),
    .S(net138),
    .X(_0525_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4320_ (.A0(rf_reg[577]),
    .A1(net329),
    .S(net138),
    .X(_0526_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4321_ (.A0(rf_reg[578]),
    .A1(net346),
    .S(net136),
    .X(_0527_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4322_ (.A0(rf_reg[579]),
    .A1(net331),
    .S(net139),
    .X(_0528_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4323_ (.A0(net333),
    .A1(rf_reg[57]),
    .S(net22),
    .X(_0529_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4324_ (.A0(rf_reg[580]),
    .A1(net337),
    .S(net137),
    .X(_0530_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4325_ (.A0(rf_reg[581]),
    .A1(net342),
    .S(net138),
    .X(_0531_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4326_ (.A0(rf_reg[582]),
    .A1(net326),
    .S(net136),
    .X(_0532_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4327_ (.A0(rf_reg[583]),
    .A1(net340),
    .S(net138),
    .X(_0533_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_109_clk_i (.X(clknet_leaf_109_clk_i),
    .A(clknet_5_16__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4329_ (.A0(rf_reg[584]),
    .A1(net341),
    .S(net136),
    .X(_0534_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_108_clk_i (.X(clknet_leaf_108_clk_i),
    .A(clknet_5_16__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4331_ (.A0(rf_reg[585]),
    .A1(net347),
    .S(net136),
    .X(_0535_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_107_clk_i (.X(clknet_leaf_107_clk_i),
    .A(clknet_5_16__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_106_clk_i (.X(clknet_leaf_106_clk_i),
    .A(clknet_5_16__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4334_ (.A0(rf_reg[586]),
    .A1(net327),
    .S(net140),
    .X(_0536_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_105_clk_i (.X(clknet_leaf_105_clk_i),
    .A(clknet_5_16__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4336_ (.A0(rf_reg[587]),
    .A1(net317),
    .S(net138),
    .X(_0537_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_104_clk_i (.X(clknet_leaf_104_clk_i),
    .A(clknet_5_17__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4338_ (.A0(rf_reg[588]),
    .A1(net322),
    .S(net140),
    .X(_0538_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_103_clk_i (.X(clknet_leaf_103_clk_i),
    .A(clknet_5_17__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4340_ (.A0(rf_reg[589]),
    .A1(net345),
    .S(net139),
    .X(_0539_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4341_ (.A0(net343),
    .A1(rf_reg[58]),
    .S(net21),
    .X(_0540_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_102_clk_i (.X(clknet_leaf_102_clk_i),
    .A(clknet_5_17__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4343_ (.A0(rf_reg[590]),
    .A1(net321),
    .S(net137),
    .X(_0541_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_101_clk_i (.X(clknet_leaf_101_clk_i),
    .A(clknet_5_20__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4345_ (.A0(rf_reg[591]),
    .A1(net332),
    .S(net137),
    .X(_0542_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_100_clk_i (.X(clknet_leaf_100_clk_i),
    .A(clknet_5_20__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4347_ (.A0(rf_reg[592]),
    .A1(net320),
    .S(net138),
    .X(_0543_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_99_clk_i (.X(clknet_leaf_99_clk_i),
    .A(clknet_5_20__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4349_ (.A0(rf_reg[593]),
    .A1(net330),
    .S(net136),
    .X(_0544_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_98_clk_i (.X(clknet_leaf_98_clk_i),
    .A(clknet_5_21__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4351_ (.A0(rf_reg[594]),
    .A1(net318),
    .S(net137),
    .X(_0545_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_97_clk_i (.X(clknet_leaf_97_clk_i),
    .A(clknet_5_21__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4353_ (.A0(rf_reg[595]),
    .A1(net325),
    .S(net138),
    .X(_0546_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_96_clk_i (.X(clknet_leaf_96_clk_i),
    .A(clknet_5_21__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_95_clk_i (.X(clknet_leaf_95_clk_i),
    .A(clknet_5_21__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4356_ (.A0(rf_reg[596]),
    .A1(net344),
    .S(net139),
    .X(_0547_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_94_clk_i (.X(clknet_leaf_94_clk_i),
    .A(clknet_5_20__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4358_ (.A0(rf_reg[597]),
    .A1(net334),
    .S(net136),
    .X(_0548_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_93_clk_i (.X(clknet_leaf_93_clk_i),
    .A(clknet_5_22__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4360_ (.A0(rf_reg[598]),
    .A1(net338),
    .S(net136),
    .X(_0549_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_92_clk_i (.X(clknet_leaf_92_clk_i),
    .A(clknet_5_22__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4362_ (.A0(rf_reg[599]),
    .A1(net324),
    .S(net139),
    .X(_0550_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4363_ (.A0(net316),
    .A1(rf_reg[59]),
    .S(net24),
    .X(_0551_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_91_clk_i (.X(clknet_leaf_91_clk_i),
    .A(clknet_5_23__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4365_ (.A0(rf_reg[600]),
    .A1(net336),
    .S(net139),
    .X(_0552_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_90_clk_i (.X(clknet_leaf_90_clk_i),
    .A(clknet_5_23__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4367_ (.A0(rf_reg[601]),
    .A1(net333),
    .S(net140),
    .X(_0553_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_89_clk_i (.X(clknet_leaf_89_clk_i),
    .A(clknet_5_23__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4369_ (.A0(rf_reg[602]),
    .A1(net343),
    .S(net137),
    .X(_0554_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_88_clk_i (.X(clknet_leaf_88_clk_i),
    .A(clknet_5_23__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4371_ (.A0(rf_reg[603]),
    .A1(net316),
    .S(net138),
    .X(_0555_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_87_clk_i (.X(clknet_leaf_87_clk_i),
    .A(clknet_5_22__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4373_ (.A0(rf_reg[604]),
    .A1(net339),
    .S(net139),
    .X(_0556_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_86_clk_i (.X(clknet_leaf_86_clk_i),
    .A(clknet_5_22__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4375_ (.A0(rf_reg[605]),
    .A1(net335),
    .S(net136),
    .X(_0557_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_85_clk_i (.X(clknet_leaf_85_clk_i),
    .A(clknet_5_19__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4377_ (.A0(rf_reg[606]),
    .A1(net319),
    .S(net137),
    .X(_0558_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_84_clk_i (.X(clknet_leaf_84_clk_i),
    .A(clknet_5_19__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4379_ (.A0(rf_reg[607]),
    .A1(net323),
    .S(net137),
    .X(_0559_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4380_ (.A(_2963_),
    .B(_3104_),
    .Y(_3133_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_83_clk_i (.X(clknet_leaf_83_clk_i),
    .A(clknet_5_19__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4382_ (.A0(rf_reg[608]),
    .A1(net328),
    .S(net133),
    .X(_0560_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4383_ (.A0(rf_reg[609]),
    .A1(net329),
    .S(net133),
    .X(_0561_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4384_ (.A0(net339),
    .A1(rf_reg[60]),
    .S(net23),
    .X(_0562_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4385_ (.A0(rf_reg[610]),
    .A1(net346),
    .S(net131),
    .X(_0563_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4386_ (.A0(rf_reg[611]),
    .A1(net331),
    .S(net134),
    .X(_0564_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_82_clk_i (.X(clknet_leaf_82_clk_i),
    .A(clknet_5_18__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4388_ (.A0(rf_reg[612]),
    .A1(net337),
    .S(net132),
    .X(_0565_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_81_clk_i (.X(clknet_leaf_81_clk_i),
    .A(clknet_5_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4390_ (.A0(rf_reg[613]),
    .A1(net342),
    .S(net134),
    .X(_0566_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_80_clk_i (.X(clknet_leaf_80_clk_i),
    .A(clknet_5_24__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4392_ (.A0(rf_reg[614]),
    .A1(net326),
    .S(net131),
    .X(_0567_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_79_clk_i (.X(clknet_leaf_79_clk_i),
    .A(clknet_5_25__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4394_ (.A0(rf_reg[615]),
    .A1(net340),
    .S(net133),
    .X(_0568_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4395_ (.A0(rf_reg[616]),
    .A1(net341),
    .S(net131),
    .X(_0569_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4396_ (.A0(rf_reg[617]),
    .A1(net347),
    .S(net131),
    .X(_0570_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_78_clk_i (.X(clknet_leaf_78_clk_i),
    .A(clknet_5_25__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4398_ (.A0(rf_reg[618]),
    .A1(net327),
    .S(net135),
    .X(_0571_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4399_ (.A0(rf_reg[619]),
    .A1(net317),
    .S(net133),
    .X(_0572_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4400_ (.A0(net335),
    .A1(rf_reg[61]),
    .S(net21),
    .X(_0573_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4401_ (.A0(rf_reg[620]),
    .A1(net322),
    .S(net132),
    .X(_0574_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4402_ (.A0(rf_reg[621]),
    .A1(net345),
    .S(net134),
    .X(_0575_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4403_ (.A0(rf_reg[622]),
    .A1(net321),
    .S(net132),
    .X(_0576_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4404_ (.A0(rf_reg[623]),
    .A1(net332),
    .S(net132),
    .X(_0577_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4405_ (.A0(rf_reg[624]),
    .A1(net320),
    .S(net133),
    .X(_0578_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4406_ (.A0(rf_reg[625]),
    .A1(net330),
    .S(net131),
    .X(_0579_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4407_ (.A0(rf_reg[626]),
    .A1(net318),
    .S(net133),
    .X(_0580_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4408_ (.A0(rf_reg[627]),
    .A1(net325),
    .S(net133),
    .X(_0581_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_77_clk_i (.X(clknet_leaf_77_clk_i),
    .A(clknet_5_25__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4410_ (.A0(rf_reg[628]),
    .A1(net344),
    .S(net134),
    .X(_0582_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4411_ (.A0(rf_reg[629]),
    .A1(net334),
    .S(net131),
    .X(_0583_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4412_ (.A0(net319),
    .A1(rf_reg[62]),
    .S(net22),
    .X(_0584_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4413_ (.A0(rf_reg[630]),
    .A1(net338),
    .S(net131),
    .X(_0585_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4414_ (.A0(rf_reg[631]),
    .A1(net324),
    .S(net134),
    .X(_0586_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4415_ (.A0(rf_reg[632]),
    .A1(net336),
    .S(net134),
    .X(_0587_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4416_ (.A0(rf_reg[633]),
    .A1(net333),
    .S(net135),
    .X(_0588_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4417_ (.A0(rf_reg[634]),
    .A1(net343),
    .S(net132),
    .X(_0589_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4418_ (.A0(rf_reg[635]),
    .A1(net316),
    .S(net133),
    .X(_0590_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4419_ (.A0(rf_reg[636]),
    .A1(net339),
    .S(net134),
    .X(_0591_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4420_ (.A0(rf_reg[637]),
    .A1(net335),
    .S(net131),
    .X(_0592_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4421_ (.A0(rf_reg[638]),
    .A1(net319),
    .S(net132),
    .X(_0593_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4422_ (.A0(rf_reg[639]),
    .A1(net323),
    .S(net132),
    .X(_0594_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4423_ (.A0(net323),
    .A1(rf_reg[63]),
    .S(net22),
    .X(_0595_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_76_clk_i (.X(clknet_leaf_76_clk_i),
    .A(clknet_5_28__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 _4425_ (.Y(_3142_),
    .B(_3018_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(_3091_));
 sg13g2_nor2_1 _4426_ (.A(_3016_),
    .B(_3142_),
    .Y(_3143_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_75_clk_i (.X(clknet_leaf_75_clk_i),
    .A(clknet_5_28__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4428_ (.A0(rf_reg[640]),
    .A1(net328),
    .S(net129),
    .X(_0596_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_74_clk_i (.X(clknet_leaf_74_clk_i),
    .A(clknet_5_28__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4430_ (.A0(rf_reg[641]),
    .A1(net329),
    .S(net129),
    .X(_0597_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_73_clk_i (.X(clknet_leaf_73_clk_i),
    .A(clknet_5_29__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4432_ (.A0(rf_reg[642]),
    .A1(net346),
    .S(net126),
    .X(_0598_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_72_clk_i (.X(clknet_leaf_72_clk_i),
    .A(clknet_5_29__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4434_ (.A0(rf_reg[643]),
    .A1(net331),
    .S(net128),
    .X(_0599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4435_ (.A0(rf_reg[644]),
    .A1(net337),
    .S(net126),
    .X(_0600_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4436_ (.A0(rf_reg[645]),
    .A1(net342),
    .S(net128),
    .X(_0601_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4437_ (.A0(rf_reg[646]),
    .A1(net326),
    .S(net127),
    .X(_0602_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4438_ (.A0(rf_reg[647]),
    .A1(net340),
    .S(net128),
    .X(_0603_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4439_ (.A0(rf_reg[648]),
    .A1(net341),
    .S(net127),
    .X(_0604_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4440_ (.A0(rf_reg[649]),
    .A1(net347),
    .S(net126),
    .X(_0605_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _4441_ (.VSS(VSS),
    .VDD(VDD),
    .X(_3148_),
    .B(_3016_),
    .A(_2967_));
 sg13g2_buf_16 clkbuf_leaf_71_clk_i (.X(clknet_leaf_71_clk_i),
    .A(clknet_5_29__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_70_clk_i (.X(clknet_leaf_70_clk_i),
    .A(clknet_5_29__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4444_ (.A0(net328),
    .A1(rf_reg[64]),
    .S(net124),
    .X(_0606_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_69_clk_i (.X(clknet_leaf_69_clk_i),
    .A(clknet_5_28__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4446_ (.A0(rf_reg[650]),
    .A1(net327),
    .S(net127),
    .X(_0607_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4447_ (.A0(rf_reg[651]),
    .A1(net317),
    .S(net129),
    .X(_0608_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4448_ (.A0(rf_reg[652]),
    .A1(net322),
    .S(net127),
    .X(_0609_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4449_ (.A0(rf_reg[653]),
    .A1(net345),
    .S(net128),
    .X(_0610_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4450_ (.A0(rf_reg[654]),
    .A1(net321),
    .S(net129),
    .X(_0611_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4451_ (.A0(rf_reg[655]),
    .A1(net332),
    .S(net129),
    .X(_0612_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4452_ (.A0(rf_reg[656]),
    .A1(net320),
    .S(net128),
    .X(_0613_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4453_ (.A0(rf_reg[657]),
    .A1(net330),
    .S(net126),
    .X(_0614_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4454_ (.A0(rf_reg[658]),
    .A1(net318),
    .S(net129),
    .X(_0615_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4455_ (.A0(rf_reg[659]),
    .A1(net325),
    .S(net129),
    .X(_0616_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4456_ (.A0(net329),
    .A1(rf_reg[65]),
    .S(net124),
    .X(_0617_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_68_clk_i (.X(clknet_leaf_68_clk_i),
    .A(clknet_5_30__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4458_ (.A0(rf_reg[660]),
    .A1(net344),
    .S(net130),
    .X(_0618_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4459_ (.A0(rf_reg[661]),
    .A1(net334),
    .S(net126),
    .X(_0619_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4460_ (.A0(rf_reg[662]),
    .A1(net338),
    .S(net126),
    .X(_0620_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4461_ (.A0(rf_reg[663]),
    .A1(net324),
    .S(net130),
    .X(_0621_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4462_ (.A0(rf_reg[664]),
    .A1(net336),
    .S(net128),
    .X(_0622_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4463_ (.A0(rf_reg[665]),
    .A1(net333),
    .S(net127),
    .X(_0623_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4464_ (.A0(rf_reg[666]),
    .A1(net343),
    .S(net126),
    .X(_0624_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4465_ (.A0(rf_reg[667]),
    .A1(net316),
    .S(net128),
    .X(_0625_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4466_ (.A0(rf_reg[668]),
    .A1(net339),
    .S(net128),
    .X(_0626_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4467_ (.A0(rf_reg[669]),
    .A1(net335),
    .S(net126),
    .X(_0627_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4468_ (.A0(net346),
    .A1(rf_reg[66]),
    .S(net121),
    .X(_0628_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4469_ (.A0(rf_reg[670]),
    .A1(net319),
    .S(net127),
    .X(_0629_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4470_ (.A0(rf_reg[671]),
    .A1(net323),
    .S(net127),
    .X(_0630_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4471_ (.A(_2963_),
    .B(_3142_),
    .Y(_3153_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_67_clk_i (.X(clknet_leaf_67_clk_i),
    .A(clknet_5_31__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4473_ (.A0(rf_reg[672]),
    .A1(net328),
    .S(net119),
    .X(_0631_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4474_ (.A0(rf_reg[673]),
    .A1(net329),
    .S(net119),
    .X(_0632_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4475_ (.A0(rf_reg[674]),
    .A1(net346),
    .S(net116),
    .X(_0633_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4476_ (.A0(rf_reg[675]),
    .A1(net331),
    .S(net118),
    .X(_0634_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4477_ (.A0(rf_reg[676]),
    .A1(net337),
    .S(net116),
    .X(_0635_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4478_ (.A0(rf_reg[677]),
    .A1(net342),
    .S(net118),
    .X(_0636_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4479_ (.A0(rf_reg[678]),
    .A1(net326),
    .S(net117),
    .X(_0637_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4480_ (.A0(rf_reg[679]),
    .A1(net340),
    .S(net118),
    .X(_0638_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4481_ (.A0(net331),
    .A1(rf_reg[67]),
    .S(net123),
    .X(_0639_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4482_ (.A0(rf_reg[680]),
    .A1(net341),
    .S(net117),
    .X(_0640_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4483_ (.A0(rf_reg[681]),
    .A1(net347),
    .S(net116),
    .X(_0641_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_66_clk_i (.X(clknet_leaf_66_clk_i),
    .A(clknet_5_31__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4485_ (.A0(rf_reg[682]),
    .A1(net327),
    .S(net117),
    .X(_0642_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4486_ (.A0(rf_reg[683]),
    .A1(net317),
    .S(net119),
    .X(_0643_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4487_ (.A0(rf_reg[684]),
    .A1(net322),
    .S(net117),
    .X(_0644_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4488_ (.A0(rf_reg[685]),
    .A1(net345),
    .S(net118),
    .X(_0645_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4489_ (.A0(rf_reg[686]),
    .A1(net321),
    .S(net119),
    .X(_0646_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4490_ (.A0(rf_reg[687]),
    .A1(net332),
    .S(net119),
    .X(_0647_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4491_ (.A0(rf_reg[688]),
    .A1(net320),
    .S(net118),
    .X(_0648_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4492_ (.A0(rf_reg[689]),
    .A1(net330),
    .S(net116),
    .X(_0649_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4493_ (.A0(net337),
    .A1(rf_reg[68]),
    .S(net121),
    .X(_0650_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4494_ (.A0(rf_reg[690]),
    .A1(net318),
    .S(net119),
    .X(_0651_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4495_ (.A0(rf_reg[691]),
    .A1(net325),
    .S(net119),
    .X(_0652_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_65_clk_i (.X(clknet_leaf_65_clk_i),
    .A(clknet_5_31__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4497_ (.A0(rf_reg[692]),
    .A1(net344),
    .S(net120),
    .X(_0653_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4498_ (.A0(rf_reg[693]),
    .A1(net334),
    .S(net116),
    .X(_0654_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4499_ (.A0(rf_reg[694]),
    .A1(net338),
    .S(net116),
    .X(_0655_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4500_ (.A0(rf_reg[695]),
    .A1(net324),
    .S(net120),
    .X(_0656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4501_ (.A0(rf_reg[696]),
    .A1(net336),
    .S(net118),
    .X(_0657_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4502_ (.A0(rf_reg[697]),
    .A1(net333),
    .S(net117),
    .X(_0658_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4503_ (.A0(rf_reg[698]),
    .A1(net343),
    .S(net116),
    .X(_0659_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4504_ (.A0(rf_reg[699]),
    .A1(net316),
    .S(net118),
    .X(_0660_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4505_ (.A0(net342),
    .A1(rf_reg[69]),
    .S(net123),
    .X(_0661_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4506_ (.A0(rf_reg[700]),
    .A1(net339),
    .S(net118),
    .X(_0662_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4507_ (.A0(rf_reg[701]),
    .A1(net335),
    .S(net116),
    .X(_0663_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4508_ (.A0(rf_reg[702]),
    .A1(net319),
    .S(net117),
    .X(_0664_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4509_ (.A0(rf_reg[703]),
    .A1(net323),
    .S(net117),
    .X(_0665_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4510_ (.A(_2950_),
    .B(_3016_),
    .Y(_3157_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_64_clk_i (.X(clknet_leaf_64_clk_i),
    .A(clknet_5_31__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4512_ (.A0(rf_reg[704]),
    .A1(net328),
    .S(net114),
    .X(_0666_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4513_ (.A0(rf_reg[705]),
    .A1(net329),
    .S(net114),
    .X(_0667_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4514_ (.A0(rf_reg[706]),
    .A1(net346),
    .S(net111),
    .X(_0668_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4515_ (.A0(rf_reg[707]),
    .A1(net331),
    .S(net113),
    .X(_0669_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4516_ (.A0(rf_reg[708]),
    .A1(net337),
    .S(net111),
    .X(_0670_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4517_ (.A0(rf_reg[709]),
    .A1(net342),
    .S(net113),
    .X(_0671_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4518_ (.A0(net326),
    .A1(rf_reg[70]),
    .S(net121),
    .X(_0672_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4519_ (.A0(rf_reg[710]),
    .A1(net326),
    .S(net112),
    .X(_0673_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4520_ (.A0(rf_reg[711]),
    .A1(net340),
    .S(net113),
    .X(_0674_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4521_ (.A0(rf_reg[712]),
    .A1(net341),
    .S(net112),
    .X(_0675_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4522_ (.A0(rf_reg[713]),
    .A1(net347),
    .S(net111),
    .X(_0676_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_63_clk_i (.X(clknet_leaf_63_clk_i),
    .A(clknet_5_30__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4524_ (.A0(rf_reg[714]),
    .A1(net327),
    .S(net114),
    .X(_0677_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4525_ (.A0(rf_reg[715]),
    .A1(net317),
    .S(net114),
    .X(_0678_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4526_ (.A0(rf_reg[716]),
    .A1(net322),
    .S(net112),
    .X(_0679_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4527_ (.A0(rf_reg[717]),
    .A1(net345),
    .S(net113),
    .X(_0680_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4528_ (.A0(rf_reg[718]),
    .A1(net321),
    .S(net114),
    .X(_0681_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4529_ (.A0(rf_reg[719]),
    .A1(net332),
    .S(net112),
    .X(_0682_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4530_ (.A0(net340),
    .A1(rf_reg[71]),
    .S(net123),
    .X(_0683_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4531_ (.A0(rf_reg[720]),
    .A1(net320),
    .S(net113),
    .X(_0684_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4532_ (.A0(rf_reg[721]),
    .A1(net330),
    .S(net111),
    .X(_0685_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4533_ (.A0(rf_reg[722]),
    .A1(net318),
    .S(net114),
    .X(_0686_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4534_ (.A0(rf_reg[723]),
    .A1(net325),
    .S(net114),
    .X(_0687_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_62_clk_i (.X(clknet_leaf_62_clk_i),
    .A(clknet_5_30__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4536_ (.A0(rf_reg[724]),
    .A1(net344),
    .S(net115),
    .X(_0688_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4537_ (.A0(rf_reg[725]),
    .A1(net334),
    .S(net111),
    .X(_0689_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4538_ (.A0(rf_reg[726]),
    .A1(net338),
    .S(net111),
    .X(_0690_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4539_ (.A0(rf_reg[727]),
    .A1(net324),
    .S(net115),
    .X(_0691_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4540_ (.A0(rf_reg[728]),
    .A1(net336),
    .S(net113),
    .X(_0692_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4541_ (.A0(rf_reg[729]),
    .A1(net333),
    .S(net112),
    .X(_0693_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4542_ (.A0(net341),
    .A1(rf_reg[72]),
    .S(net121),
    .X(_0694_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4543_ (.A0(rf_reg[730]),
    .A1(net343),
    .S(net111),
    .X(_0695_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4544_ (.A0(rf_reg[731]),
    .A1(net316),
    .S(net113),
    .X(_0696_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4545_ (.A0(rf_reg[732]),
    .A1(net339),
    .S(net113),
    .X(_0697_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4546_ (.A0(rf_reg[733]),
    .A1(net335),
    .S(net111),
    .X(_0698_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4547_ (.A0(rf_reg[734]),
    .A1(net319),
    .S(net112),
    .X(_0699_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4548_ (.A0(rf_reg[735]),
    .A1(net323),
    .S(net112),
    .X(_0700_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4549_ (.A(_2950_),
    .B(_2963_),
    .Y(_3161_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_61_clk_i (.X(clknet_leaf_61_clk_i),
    .A(clknet_5_30__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4551_ (.A0(rf_reg[736]),
    .A1(net328),
    .S(net109),
    .X(_0701_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4552_ (.A0(rf_reg[737]),
    .A1(net329),
    .S(net109),
    .X(_0702_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4553_ (.A0(rf_reg[738]),
    .A1(net346),
    .S(net106),
    .X(_0703_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4554_ (.A0(rf_reg[739]),
    .A1(net331),
    .S(net108),
    .X(_0704_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4555_ (.A0(net347),
    .A1(rf_reg[73]),
    .S(net121),
    .X(_0705_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4556_ (.A0(rf_reg[740]),
    .A1(net337),
    .S(net106),
    .X(_0706_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4557_ (.A0(rf_reg[741]),
    .A1(net342),
    .S(net108),
    .X(_0707_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4558_ (.A0(rf_reg[742]),
    .A1(net326),
    .S(net107),
    .X(_0708_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4559_ (.A0(rf_reg[743]),
    .A1(net340),
    .S(net108),
    .X(_0709_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4560_ (.A0(rf_reg[744]),
    .A1(net341),
    .S(net107),
    .X(_0710_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4561_ (.A0(rf_reg[745]),
    .A1(net347),
    .S(net106),
    .X(_0711_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_60_clk_i (.X(clknet_leaf_60_clk_i),
    .A(clknet_5_27__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4563_ (.A0(rf_reg[746]),
    .A1(net327),
    .S(net107),
    .X(_0712_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4564_ (.A0(rf_reg[747]),
    .A1(net317),
    .S(net109),
    .X(_0713_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4565_ (.A0(rf_reg[748]),
    .A1(net322),
    .S(net107),
    .X(_0714_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4566_ (.A0(rf_reg[749]),
    .A1(net345),
    .S(net108),
    .X(_0715_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_59_clk_i (.X(clknet_leaf_59_clk_i),
    .A(clknet_5_27__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4568_ (.A0(net327),
    .A1(rf_reg[74]),
    .S(net122),
    .X(_0716_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4569_ (.A0(rf_reg[750]),
    .A1(net321),
    .S(net109),
    .X(_0717_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4570_ (.A0(rf_reg[751]),
    .A1(net332),
    .S(net107),
    .X(_0718_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4571_ (.A0(rf_reg[752]),
    .A1(net320),
    .S(net108),
    .X(_0719_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4572_ (.A0(rf_reg[753]),
    .A1(net330),
    .S(net106),
    .X(_0720_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4573_ (.A0(rf_reg[754]),
    .A1(net318),
    .S(net109),
    .X(_0721_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4574_ (.A0(rf_reg[755]),
    .A1(net325),
    .S(net109),
    .X(_0722_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_58_clk_i (.X(clknet_leaf_58_clk_i),
    .A(clknet_5_27__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4576_ (.A0(rf_reg[756]),
    .A1(net344),
    .S(net109),
    .X(_0723_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4577_ (.A0(rf_reg[757]),
    .A1(net334),
    .S(net106),
    .X(_0724_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4578_ (.A0(rf_reg[758]),
    .A1(net338),
    .S(net106),
    .X(_0725_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4579_ (.A0(rf_reg[759]),
    .A1(net324),
    .S(net110),
    .X(_0726_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4580_ (.A0(net317),
    .A1(rf_reg[75]),
    .S(net124),
    .X(_0727_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4581_ (.A0(rf_reg[760]),
    .A1(net336),
    .S(net108),
    .X(_0728_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4582_ (.A0(rf_reg[761]),
    .A1(net333),
    .S(net107),
    .X(_0729_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4583_ (.A0(rf_reg[762]),
    .A1(net343),
    .S(net106),
    .X(_0730_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4584_ (.A0(rf_reg[763]),
    .A1(net316),
    .S(net108),
    .X(_0731_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4585_ (.A0(rf_reg[764]),
    .A1(net339),
    .S(net108),
    .X(_0732_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4586_ (.A0(rf_reg[765]),
    .A1(net335),
    .S(net106),
    .X(_0733_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4587_ (.A0(rf_reg[766]),
    .A1(net319),
    .S(net107),
    .X(_0734_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4588_ (.A0(rf_reg[767]),
    .A1(net323),
    .S(net107),
    .X(_0735_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _4589_ (.Y(_3166_),
    .B(_3092_),
    .A_N(_3049_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_57_clk_i (.X(clknet_leaf_57_clk_i),
    .A(clknet_5_26__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_56_clk_i (.X(clknet_leaf_56_clk_i),
    .A(clknet_5_26__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4592_ (.A0(net328),
    .A1(rf_reg[768]),
    .S(net104),
    .X(_0736_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4593_ (.A0(net329),
    .A1(rf_reg[769]),
    .S(net104),
    .X(_0737_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4594_ (.A0(net322),
    .A1(rf_reg[76]),
    .S(net122),
    .X(_0738_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4595_ (.A0(net346),
    .A1(rf_reg[770]),
    .S(net101),
    .X(_0739_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4596_ (.A0(net331),
    .A1(rf_reg[771]),
    .S(net103),
    .X(_0740_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4597_ (.A0(net337),
    .A1(rf_reg[772]),
    .S(net101),
    .X(_0741_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4598_ (.A0(net342),
    .A1(rf_reg[773]),
    .S(net103),
    .X(_0742_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4599_ (.A0(net326),
    .A1(rf_reg[774]),
    .S(net101),
    .X(_0743_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4600_ (.A0(net340),
    .A1(rf_reg[775]),
    .S(net103),
    .X(_0744_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4601_ (.A0(net341),
    .A1(rf_reg[776]),
    .S(net101),
    .X(_0745_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4602_ (.A0(net347),
    .A1(rf_reg[777]),
    .S(net101),
    .X(_0746_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_55_clk_i (.X(clknet_leaf_55_clk_i),
    .A(clknet_5_26__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4604_ (.A0(net327),
    .A1(rf_reg[778]),
    .S(net102),
    .X(_0747_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4605_ (.A0(net317),
    .A1(rf_reg[779]),
    .S(net104),
    .X(_0748_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4606_ (.A0(net345),
    .A1(rf_reg[77]),
    .S(net123),
    .X(_0749_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4607_ (.A0(net322),
    .A1(rf_reg[780]),
    .S(net102),
    .X(_0750_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4608_ (.A0(net345),
    .A1(rf_reg[781]),
    .S(net103),
    .X(_0751_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4609_ (.A0(net321),
    .A1(rf_reg[782]),
    .S(net104),
    .X(_0752_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4610_ (.A0(net332),
    .A1(rf_reg[783]),
    .S(net102),
    .X(_0753_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4611_ (.A0(net320),
    .A1(rf_reg[784]),
    .S(net103),
    .X(_0754_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4612_ (.A0(net330),
    .A1(rf_reg[785]),
    .S(net102),
    .X(_0755_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4613_ (.A0(net318),
    .A1(rf_reg[786]),
    .S(net104),
    .X(_0756_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4614_ (.A0(net325),
    .A1(rf_reg[787]),
    .S(net104),
    .X(_0757_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_54_clk_i (.X(clknet_leaf_54_clk_i),
    .A(clknet_5_26__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4616_ (.A0(net344),
    .A1(rf_reg[788]),
    .S(net103),
    .X(_0758_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4617_ (.A0(net334),
    .A1(rf_reg[789]),
    .S(net102),
    .X(_0759_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4618_ (.A0(net321),
    .A1(rf_reg[78]),
    .S(net124),
    .X(_0760_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4619_ (.A0(net338),
    .A1(rf_reg[790]),
    .S(net102),
    .X(_0761_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4620_ (.A0(net324),
    .A1(rf_reg[791]),
    .S(net104),
    .X(_0762_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4621_ (.A0(net336),
    .A1(rf_reg[792]),
    .S(net105),
    .X(_0763_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4622_ (.A0(net333),
    .A1(rf_reg[793]),
    .S(net105),
    .X(_0764_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4623_ (.A0(net343),
    .A1(rf_reg[794]),
    .S(net101),
    .X(_0765_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4624_ (.A0(net316),
    .A1(rf_reg[795]),
    .S(net103),
    .X(_0766_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4625_ (.A0(net339),
    .A1(rf_reg[796]),
    .S(net103),
    .X(_0767_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4626_ (.A0(net335),
    .A1(rf_reg[797]),
    .S(net101),
    .X(_0768_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4627_ (.A0(net319),
    .A1(rf_reg[798]),
    .S(net102),
    .X(_0769_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4628_ (.A0(net323),
    .A1(rf_reg[799]),
    .S(net101),
    .X(_0770_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4629_ (.A0(net332),
    .A1(rf_reg[79]),
    .S(net124),
    .X(_0771_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _4630_ (.Y(_3171_),
    .B(_3092_),
    .A_N(_2949_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_53_clk_i (.X(clknet_leaf_53_clk_i),
    .A(clknet_5_27__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_52_clk_i (.X(clknet_leaf_52_clk_i),
    .A(clknet_5_25__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4633_ (.A0(net328),
    .A1(rf_reg[800]),
    .S(net99),
    .X(_0772_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4634_ (.A0(net329),
    .A1(rf_reg[801]),
    .S(net99),
    .X(_0773_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4635_ (.A0(net346),
    .A1(rf_reg[802]),
    .S(net96),
    .X(_0774_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4636_ (.A0(net331),
    .A1(rf_reg[803]),
    .S(net98),
    .X(_0775_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4637_ (.A0(net337),
    .A1(rf_reg[804]),
    .S(net96),
    .X(_0776_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4638_ (.A0(net342),
    .A1(rf_reg[805]),
    .S(net98),
    .X(_0777_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4639_ (.A0(net326),
    .A1(rf_reg[806]),
    .S(net96),
    .X(_0778_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4640_ (.A0(net340),
    .A1(rf_reg[807]),
    .S(net98),
    .X(_0779_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4641_ (.A0(net341),
    .A1(rf_reg[808]),
    .S(net96),
    .X(_0780_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4642_ (.A0(net347),
    .A1(rf_reg[809]),
    .S(net96),
    .X(_0781_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4643_ (.A0(net320),
    .A1(rf_reg[80]),
    .S(net123),
    .X(_0782_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_51_clk_i (.X(clknet_leaf_51_clk_i),
    .A(clknet_5_24__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4645_ (.A0(net327),
    .A1(rf_reg[810]),
    .S(net97),
    .X(_0783_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4646_ (.A0(net317),
    .A1(rf_reg[811]),
    .S(net99),
    .X(_0784_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4647_ (.A0(net322),
    .A1(rf_reg[812]),
    .S(net97),
    .X(_0785_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4648_ (.A0(net345),
    .A1(rf_reg[813]),
    .S(net98),
    .X(_0786_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4649_ (.A0(net321),
    .A1(rf_reg[814]),
    .S(net99),
    .X(_0787_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4650_ (.A0(net332),
    .A1(rf_reg[815]),
    .S(net97),
    .X(_0788_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4651_ (.A0(net320),
    .A1(rf_reg[816]),
    .S(net98),
    .X(_0789_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4652_ (.A0(net330),
    .A1(rf_reg[817]),
    .S(net97),
    .X(_0790_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4653_ (.A0(net318),
    .A1(rf_reg[818]),
    .S(net99),
    .X(_0791_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4654_ (.A0(net325),
    .A1(rf_reg[819]),
    .S(net99),
    .X(_0792_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4655_ (.A0(net330),
    .A1(rf_reg[81]),
    .S(net121),
    .X(_0793_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_50_clk_i (.X(clknet_leaf_50_clk_i),
    .A(clknet_5_24__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4657_ (.A0(net344),
    .A1(rf_reg[820]),
    .S(net98),
    .X(_0794_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4658_ (.A0(net334),
    .A1(rf_reg[821]),
    .S(net97),
    .X(_0795_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4659_ (.A0(net338),
    .A1(rf_reg[822]),
    .S(net97),
    .X(_0796_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4660_ (.A0(net324),
    .A1(rf_reg[823]),
    .S(net99),
    .X(_0797_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4661_ (.A0(net336),
    .A1(rf_reg[824]),
    .S(net100),
    .X(_0798_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4662_ (.A0(net333),
    .A1(rf_reg[825]),
    .S(net100),
    .X(_0799_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4663_ (.A0(net343),
    .A1(rf_reg[826]),
    .S(net96),
    .X(_0800_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4664_ (.A0(net316),
    .A1(rf_reg[827]),
    .S(net98),
    .X(_0801_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4665_ (.A0(net339),
    .A1(rf_reg[828]),
    .S(net98),
    .X(_0802_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4666_ (.A0(net335),
    .A1(rf_reg[829]),
    .S(net96),
    .X(_0803_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4667_ (.A0(net318),
    .A1(rf_reg[82]),
    .S(net124),
    .X(_0804_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4668_ (.A0(net319),
    .A1(rf_reg[830]),
    .S(net97),
    .X(_0805_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4669_ (.A0(net323),
    .A1(rf_reg[831]),
    .S(net96),
    .X(_0806_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4670_ (.A(_3049_),
    .B(_3104_),
    .Y(_3176_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_49_clk_i (.X(clknet_leaf_49_clk_i),
    .A(clknet_5_24__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4672_ (.A0(rf_reg[832]),
    .A1(net328),
    .S(net94),
    .X(_0807_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4673_ (.A0(rf_reg[833]),
    .A1(net329),
    .S(net94),
    .X(_0808_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4674_ (.A0(rf_reg[834]),
    .A1(net346),
    .S(net91),
    .X(_0809_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4675_ (.A0(rf_reg[835]),
    .A1(net331),
    .S(net93),
    .X(_0810_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4676_ (.A0(rf_reg[836]),
    .A1(net337),
    .S(net91),
    .X(_0811_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4677_ (.A0(rf_reg[837]),
    .A1(net342),
    .S(net93),
    .X(_0812_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4678_ (.A0(rf_reg[838]),
    .A1(net326),
    .S(net91),
    .X(_0813_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4679_ (.A0(rf_reg[839]),
    .A1(net340),
    .S(net93),
    .X(_0814_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4680_ (.A0(net325),
    .A1(rf_reg[83]),
    .S(net124),
    .X(_0815_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4681_ (.A0(rf_reg[840]),
    .A1(net341),
    .S(net91),
    .X(_0816_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4682_ (.A0(rf_reg[841]),
    .A1(net347),
    .S(net91),
    .X(_0817_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_48_clk_i (.X(clknet_leaf_48_clk_i),
    .A(clknet_5_13__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4684_ (.A0(rf_reg[842]),
    .A1(net327),
    .S(net92),
    .X(_0818_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4685_ (.A0(rf_reg[843]),
    .A1(net317),
    .S(net94),
    .X(_0819_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4686_ (.A0(rf_reg[844]),
    .A1(net322),
    .S(net92),
    .X(_0820_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4687_ (.A0(rf_reg[845]),
    .A1(net345),
    .S(net93),
    .X(_0821_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4688_ (.A0(rf_reg[846]),
    .A1(net321),
    .S(net94),
    .X(_0822_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4689_ (.A0(rf_reg[847]),
    .A1(net332),
    .S(net94),
    .X(_0823_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4690_ (.A0(rf_reg[848]),
    .A1(net320),
    .S(net93),
    .X(_0824_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4691_ (.A0(rf_reg[849]),
    .A1(net330),
    .S(net91),
    .X(_0825_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_47_clk_i (.X(clknet_leaf_47_clk_i),
    .A(clknet_5_12__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4693_ (.A0(net344),
    .A1(rf_reg[84]),
    .S(net123),
    .X(_0826_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4694_ (.A0(rf_reg[850]),
    .A1(net318),
    .S(net94),
    .X(_0827_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4695_ (.A0(rf_reg[851]),
    .A1(net325),
    .S(net94),
    .X(_0828_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_46_clk_i (.X(clknet_leaf_46_clk_i),
    .A(clknet_5_13__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4697_ (.A0(rf_reg[852]),
    .A1(net344),
    .S(net93),
    .X(_0829_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4698_ (.A0(rf_reg[853]),
    .A1(net334),
    .S(net92),
    .X(_0830_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4699_ (.A0(rf_reg[854]),
    .A1(net338),
    .S(net92),
    .X(_0831_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4700_ (.A0(rf_reg[855]),
    .A1(net324),
    .S(net95),
    .X(_0832_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4701_ (.A0(rf_reg[856]),
    .A1(net336),
    .S(net95),
    .X(_0833_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4702_ (.A0(rf_reg[857]),
    .A1(net333),
    .S(net92),
    .X(_0834_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4703_ (.A0(rf_reg[858]),
    .A1(net343),
    .S(net91),
    .X(_0835_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4704_ (.A0(rf_reg[859]),
    .A1(net316),
    .S(net93),
    .X(_0836_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4705_ (.A0(net334),
    .A1(rf_reg[85]),
    .S(net122),
    .X(_0837_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4706_ (.A0(rf_reg[860]),
    .A1(net339),
    .S(net93),
    .X(_0838_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4707_ (.A0(rf_reg[861]),
    .A1(net335),
    .S(net91),
    .X(_0839_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4708_ (.A0(rf_reg[862]),
    .A1(net319),
    .S(net92),
    .X(_0840_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4709_ (.A0(rf_reg[863]),
    .A1(net323),
    .S(net92),
    .X(_0841_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4710_ (.A(_2949_),
    .B(_3104_),
    .Y(_3181_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_45_clk_i (.X(clknet_leaf_45_clk_i),
    .A(clknet_5_13__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4712_ (.A0(rf_reg[864]),
    .A1(net328),
    .S(net89),
    .X(_0842_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4713_ (.A0(rf_reg[865]),
    .A1(net329),
    .S(net89),
    .X(_0843_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4714_ (.A0(rf_reg[866]),
    .A1(net346),
    .S(net86),
    .X(_0844_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4715_ (.A0(rf_reg[867]),
    .A1(net331),
    .S(net88),
    .X(_0845_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4716_ (.A0(rf_reg[868]),
    .A1(net337),
    .S(net86),
    .X(_0846_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4717_ (.A0(rf_reg[869]),
    .A1(net342),
    .S(net88),
    .X(_0847_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4718_ (.A0(net338),
    .A1(rf_reg[86]),
    .S(net122),
    .X(_0848_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4719_ (.A0(rf_reg[870]),
    .A1(net326),
    .S(net86),
    .X(_0849_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4720_ (.A0(rf_reg[871]),
    .A1(net340),
    .S(net88),
    .X(_0850_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4721_ (.A0(rf_reg[872]),
    .A1(net341),
    .S(net86),
    .X(_0851_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4722_ (.A0(rf_reg[873]),
    .A1(net347),
    .S(net86),
    .X(_0852_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_44_clk_i (.X(clknet_leaf_44_clk_i),
    .A(clknet_5_14__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4724_ (.A0(rf_reg[874]),
    .A1(net327),
    .S(net87),
    .X(_0853_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4725_ (.A0(rf_reg[875]),
    .A1(net317),
    .S(net89),
    .X(_0854_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4726_ (.A0(rf_reg[876]),
    .A1(net322),
    .S(net87),
    .X(_0855_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4727_ (.A0(rf_reg[877]),
    .A1(net345),
    .S(net88),
    .X(_0856_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4728_ (.A0(rf_reg[878]),
    .A1(net321),
    .S(net89),
    .X(_0857_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4729_ (.A0(rf_reg[879]),
    .A1(net332),
    .S(net89),
    .X(_0858_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4730_ (.A0(net324),
    .A1(rf_reg[87]),
    .S(net125),
    .X(_0859_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4731_ (.A0(rf_reg[880]),
    .A1(net320),
    .S(net88),
    .X(_0860_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4732_ (.A0(rf_reg[881]),
    .A1(net330),
    .S(net87),
    .X(_0861_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4733_ (.A0(rf_reg[882]),
    .A1(net318),
    .S(net89),
    .X(_0862_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4734_ (.A0(rf_reg[883]),
    .A1(net325),
    .S(net89),
    .X(_0863_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_43_clk_i (.X(clknet_leaf_43_clk_i),
    .A(clknet_5_15__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4736_ (.A0(rf_reg[884]),
    .A1(net344),
    .S(net88),
    .X(_0864_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4737_ (.A0(rf_reg[885]),
    .A1(net334),
    .S(net87),
    .X(_0865_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4738_ (.A0(rf_reg[886]),
    .A1(net338),
    .S(net87),
    .X(_0866_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4739_ (.A0(rf_reg[887]),
    .A1(net324),
    .S(net90),
    .X(_0867_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4740_ (.A0(rf_reg[888]),
    .A1(net336),
    .S(net90),
    .X(_0868_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4741_ (.A0(rf_reg[889]),
    .A1(net333),
    .S(net87),
    .X(_0869_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4742_ (.A0(net336),
    .A1(rf_reg[88]),
    .S(net125),
    .X(_0870_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4743_ (.A0(rf_reg[890]),
    .A1(net343),
    .S(net86),
    .X(_0871_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4744_ (.A0(rf_reg[891]),
    .A1(net316),
    .S(net88),
    .X(_0872_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4745_ (.A0(rf_reg[892]),
    .A1(net339),
    .S(net88),
    .X(_0873_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4746_ (.A0(rf_reg[893]),
    .A1(net335),
    .S(net86),
    .X(_0874_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4747_ (.A0(rf_reg[894]),
    .A1(net319),
    .S(net87),
    .X(_0875_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4748_ (.A0(rf_reg[895]),
    .A1(net323),
    .S(net86),
    .X(_0876_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4749_ (.A(_3049_),
    .B(_3142_),
    .Y(_3185_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_42_clk_i (.X(clknet_leaf_42_clk_i),
    .A(clknet_5_15__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4751_ (.A0(rf_reg[896]),
    .A1(net328),
    .S(net84),
    .X(_0877_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4752_ (.A0(rf_reg[897]),
    .A1(net329),
    .S(net84),
    .X(_0878_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4753_ (.A0(rf_reg[898]),
    .A1(net346),
    .S(net81),
    .X(_0879_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4754_ (.A0(rf_reg[899]),
    .A1(net331),
    .S(net83),
    .X(_0880_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4755_ (.A0(net333),
    .A1(rf_reg[89]),
    .S(net122),
    .X(_0881_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4756_ (.A0(rf_reg[900]),
    .A1(net337),
    .S(net81),
    .X(_0882_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4757_ (.A0(rf_reg[901]),
    .A1(net342),
    .S(net83),
    .X(_0883_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4758_ (.A0(rf_reg[902]),
    .A1(net326),
    .S(net81),
    .X(_0884_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4759_ (.A0(rf_reg[903]),
    .A1(net340),
    .S(net83),
    .X(_0885_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4760_ (.A0(rf_reg[904]),
    .A1(net341),
    .S(net81),
    .X(_0886_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4761_ (.A0(rf_reg[905]),
    .A1(net347),
    .S(net81),
    .X(_0887_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_41_clk_i (.X(clknet_leaf_41_clk_i),
    .A(clknet_5_15__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4763_ (.A0(rf_reg[906]),
    .A1(net327),
    .S(net82),
    .X(_0888_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4764_ (.A0(rf_reg[907]),
    .A1(net317),
    .S(net84),
    .X(_0889_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4765_ (.A0(rf_reg[908]),
    .A1(net322),
    .S(net82),
    .X(_0890_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4766_ (.A0(rf_reg[909]),
    .A1(net345),
    .S(net83),
    .X(_0891_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4767_ (.A0(net343),
    .A1(rf_reg[90]),
    .S(net122),
    .X(_0892_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4768_ (.A0(rf_reg[910]),
    .A1(net321),
    .S(net84),
    .X(_0893_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4769_ (.A0(rf_reg[911]),
    .A1(net332),
    .S(net82),
    .X(_0894_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4770_ (.A0(rf_reg[912]),
    .A1(net320),
    .S(net83),
    .X(_0895_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4771_ (.A0(rf_reg[913]),
    .A1(net330),
    .S(net81),
    .X(_0896_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4772_ (.A0(rf_reg[914]),
    .A1(net318),
    .S(net84),
    .X(_0897_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4773_ (.A0(rf_reg[915]),
    .A1(net325),
    .S(net85),
    .X(_0898_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_40_clk_i (.X(clknet_leaf_40_clk_i),
    .A(clknet_5_15__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4775_ (.A0(rf_reg[916]),
    .A1(net344),
    .S(net83),
    .X(_0899_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4776_ (.A0(rf_reg[917]),
    .A1(net334),
    .S(net82),
    .X(_0900_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4777_ (.A0(rf_reg[918]),
    .A1(net338),
    .S(net82),
    .X(_0901_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4778_ (.A0(rf_reg[919]),
    .A1(net324),
    .S(net84),
    .X(_0902_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4779_ (.A0(net316),
    .A1(rf_reg[91]),
    .S(net123),
    .X(_0903_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4780_ (.A0(rf_reg[920]),
    .A1(net336),
    .S(net83),
    .X(_0904_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4781_ (.A0(rf_reg[921]),
    .A1(net333),
    .S(net85),
    .X(_0905_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4782_ (.A0(rf_reg[922]),
    .A1(net343),
    .S(net81),
    .X(_0906_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4783_ (.A0(rf_reg[923]),
    .A1(net316),
    .S(net84),
    .X(_0907_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4784_ (.A0(rf_reg[924]),
    .A1(net339),
    .S(net83),
    .X(_0908_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4785_ (.A0(rf_reg[925]),
    .A1(net335),
    .S(net81),
    .X(_0909_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4786_ (.A0(rf_reg[926]),
    .A1(net319),
    .S(net82),
    .X(_0910_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4787_ (.A0(rf_reg[927]),
    .A1(net323),
    .S(net82),
    .X(_0911_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4788_ (.A(_2949_),
    .B(_3142_),
    .Y(_3189_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_39_clk_i (.X(clknet_leaf_39_clk_i),
    .A(clknet_5_14__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4790_ (.A0(rf_reg[928]),
    .A1(net328),
    .S(net79),
    .X(_0912_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4791_ (.A0(rf_reg[929]),
    .A1(net329),
    .S(net79),
    .X(_0913_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4792_ (.A0(net339),
    .A1(rf_reg[92]),
    .S(net123),
    .X(_0914_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4793_ (.A0(rf_reg[930]),
    .A1(net346),
    .S(net76),
    .X(_0915_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4794_ (.A0(rf_reg[931]),
    .A1(net331),
    .S(net78),
    .X(_0916_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4795_ (.A0(rf_reg[932]),
    .A1(net337),
    .S(net76),
    .X(_0917_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4796_ (.A0(rf_reg[933]),
    .A1(net342),
    .S(net78),
    .X(_0918_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4797_ (.A0(rf_reg[934]),
    .A1(net326),
    .S(net76),
    .X(_0919_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4798_ (.A0(rf_reg[935]),
    .A1(net340),
    .S(net78),
    .X(_0920_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4799_ (.A0(rf_reg[936]),
    .A1(net341),
    .S(net76),
    .X(_0921_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4800_ (.A0(rf_reg[937]),
    .A1(net347),
    .S(net76),
    .X(_0922_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_38_clk_i (.X(clknet_leaf_38_clk_i),
    .A(clknet_5_14__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4802_ (.A0(rf_reg[938]),
    .A1(net327),
    .S(net77),
    .X(_0923_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4803_ (.A0(rf_reg[939]),
    .A1(net317),
    .S(net79),
    .X(_0924_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4804_ (.A0(net335),
    .A1(rf_reg[93]),
    .S(net121),
    .X(_0925_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4805_ (.A0(rf_reg[940]),
    .A1(net322),
    .S(net77),
    .X(_0926_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4806_ (.A0(rf_reg[941]),
    .A1(net345),
    .S(net78),
    .X(_0927_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4807_ (.A0(rf_reg[942]),
    .A1(net321),
    .S(net79),
    .X(_0928_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4808_ (.A0(rf_reg[943]),
    .A1(net332),
    .S(net79),
    .X(_0929_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4809_ (.A0(rf_reg[944]),
    .A1(net320),
    .S(net78),
    .X(_0930_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4810_ (.A0(rf_reg[945]),
    .A1(net330),
    .S(net76),
    .X(_0931_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4811_ (.A0(rf_reg[946]),
    .A1(net318),
    .S(net79),
    .X(_0932_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4812_ (.A0(rf_reg[947]),
    .A1(net325),
    .S(net80),
    .X(_0933_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_37_clk_i (.X(clknet_leaf_37_clk_i),
    .A(clknet_5_14__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4814_ (.A0(rf_reg[948]),
    .A1(net344),
    .S(net78),
    .X(_0934_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4815_ (.A0(rf_reg[949]),
    .A1(net334),
    .S(net77),
    .X(_0935_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4816_ (.A0(net319),
    .A1(rf_reg[94]),
    .S(net122),
    .X(_0936_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4817_ (.A0(rf_reg[950]),
    .A1(net338),
    .S(net77),
    .X(_0937_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4818_ (.A0(rf_reg[951]),
    .A1(net324),
    .S(net79),
    .X(_0938_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4819_ (.A0(rf_reg[952]),
    .A1(net336),
    .S(net78),
    .X(_0939_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4820_ (.A0(rf_reg[953]),
    .A1(net333),
    .S(net77),
    .X(_0940_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4821_ (.A0(rf_reg[954]),
    .A1(net343),
    .S(net76),
    .X(_0941_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4822_ (.A0(rf_reg[955]),
    .A1(net316),
    .S(net80),
    .X(_0942_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4823_ (.A0(rf_reg[956]),
    .A1(net339),
    .S(net78),
    .X(_0943_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4824_ (.A0(rf_reg[957]),
    .A1(net335),
    .S(net76),
    .X(_0944_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4825_ (.A0(rf_reg[958]),
    .A1(net319),
    .S(net77),
    .X(_0945_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4826_ (.A0(rf_reg[959]),
    .A1(net323),
    .S(net77),
    .X(_0946_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4827_ (.A0(net323),
    .A1(rf_reg[95]),
    .S(net121),
    .X(_0947_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _4828_ (.A(_2950_),
    .B(_3049_),
    .Y(_3193_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_36_clk_i (.X(clknet_leaf_36_clk_i),
    .A(clknet_5_11__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4830_ (.A0(rf_reg[960]),
    .A1(net328),
    .S(net75),
    .X(_0948_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4831_ (.A0(rf_reg[961]),
    .A1(net329),
    .S(net75),
    .X(_0949_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4832_ (.A0(rf_reg[962]),
    .A1(net346),
    .S(net71),
    .X(_0950_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4833_ (.A0(rf_reg[963]),
    .A1(net331),
    .S(net74),
    .X(_0951_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4834_ (.A0(rf_reg[964]),
    .A1(net337),
    .S(net72),
    .X(_0952_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4835_ (.A0(rf_reg[965]),
    .A1(net342),
    .S(net74),
    .X(_0953_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4836_ (.A0(rf_reg[966]),
    .A1(net326),
    .S(net72),
    .X(_0954_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4837_ (.A0(rf_reg[967]),
    .A1(net340),
    .S(net74),
    .X(_0955_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4838_ (.A0(rf_reg[968]),
    .A1(net341),
    .S(net71),
    .X(_0956_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4839_ (.A0(rf_reg[969]),
    .A1(net347),
    .S(net71),
    .X(_0957_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4840_ (.A0(rf_reg[96]),
    .A1(net328),
    .S(net64),
    .X(_0958_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_35_clk_i (.X(clknet_leaf_35_clk_i),
    .A(clknet_5_11__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4842_ (.A0(rf_reg[970]),
    .A1(net327),
    .S(net73),
    .X(_0959_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4843_ (.A0(rf_reg[971]),
    .A1(net317),
    .S(net75),
    .X(_0960_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4844_ (.A0(rf_reg[972]),
    .A1(net322),
    .S(net71),
    .X(_0961_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4845_ (.A0(rf_reg[973]),
    .A1(net345),
    .S(net74),
    .X(_0962_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4846_ (.A0(rf_reg[974]),
    .A1(net321),
    .S(net73),
    .X(_0963_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4847_ (.A0(rf_reg[975]),
    .A1(net332),
    .S(net73),
    .X(_0964_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4848_ (.A0(rf_reg[976]),
    .A1(net320),
    .S(net74),
    .X(_0965_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4849_ (.A0(rf_reg[977]),
    .A1(net330),
    .S(net72),
    .X(_0966_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4850_ (.A0(rf_reg[978]),
    .A1(net318),
    .S(net75),
    .X(_0967_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4851_ (.A0(rf_reg[979]),
    .A1(net325),
    .S(net75),
    .X(_0968_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4852_ (.A0(rf_reg[97]),
    .A1(net329),
    .S(net64),
    .X(_0969_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_34_clk_i (.X(clknet_leaf_34_clk_i),
    .A(clknet_5_10__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4854_ (.A0(rf_reg[980]),
    .A1(net344),
    .S(net74),
    .X(_0970_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4855_ (.A0(rf_reg[981]),
    .A1(net334),
    .S(net72),
    .X(_0971_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4856_ (.A0(rf_reg[982]),
    .A1(net338),
    .S(net72),
    .X(_0972_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4857_ (.A0(rf_reg[983]),
    .A1(net324),
    .S(net75),
    .X(_0973_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4858_ (.A0(rf_reg[984]),
    .A1(net336),
    .S(net74),
    .X(_0974_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4859_ (.A0(rf_reg[985]),
    .A1(net333),
    .S(net73),
    .X(_0975_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4860_ (.A0(rf_reg[986]),
    .A1(net343),
    .S(net71),
    .X(_0976_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4861_ (.A0(rf_reg[987]),
    .A1(net316),
    .S(net75),
    .X(_0977_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4862_ (.A0(rf_reg[988]),
    .A1(net339),
    .S(net74),
    .X(_0978_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4863_ (.A0(rf_reg[989]),
    .A1(net335),
    .S(net71),
    .X(_0979_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4864_ (.A0(rf_reg[98]),
    .A1(net346),
    .S(net61),
    .X(_0980_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4865_ (.A0(rf_reg[990]),
    .A1(net319),
    .S(net71),
    .X(_0981_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4866_ (.A0(rf_reg[991]),
    .A1(net323),
    .S(net71),
    .X(_0982_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4867_ (.A0(rf_reg[992]),
    .A1(net328),
    .S(net160),
    .X(_0983_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4868_ (.A0(rf_reg[993]),
    .A1(net329),
    .S(net160),
    .X(_0984_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4869_ (.A0(rf_reg[994]),
    .A1(net346),
    .S(net156),
    .X(_0985_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4870_ (.A0(rf_reg[995]),
    .A1(net331),
    .S(net160),
    .X(_0986_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4871_ (.A0(rf_reg[996]),
    .A1(net337),
    .S(net157),
    .X(_0987_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4872_ (.A0(rf_reg[997]),
    .A1(net342),
    .S(net159),
    .X(_0988_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4873_ (.A0(rf_reg[998]),
    .A1(net326),
    .S(net156),
    .X(_0989_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4874_ (.A0(rf_reg[999]),
    .A1(net340),
    .S(net159),
    .X(_0990_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4875_ (.A0(rf_reg[99]),
    .A1(net331),
    .S(net63),
    .X(_0991_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_33_clk_i (.X(clknet_leaf_33_clk_i),
    .A(clknet_5_10__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _4877_ (.A(raddr_a_i[1]),
    .B(raddr_a_i[2]),
    .X(_0993_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_32_clk_i (.X(clknet_leaf_32_clk_i),
    .A(clknet_5_10__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_31_clk_i (.X(clknet_leaf_31_clk_i),
    .A(clknet_5_10__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_30_clk_i (.X(clknet_leaf_30_clk_i),
    .A(clknet_5_11__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_29_clk_i (.X(clknet_leaf_29_clk_i),
    .A(clknet_5_11__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_28_clk_i (.X(clknet_leaf_28_clk_i),
    .A(clknet_5_8__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_27_clk_i (.X(clknet_leaf_27_clk_i),
    .A(clknet_5_8__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4884_ (.A0(rf_reg[479]),
    .A1(rf_reg[511]),
    .S(raddr_a_i[0]),
    .X(_1000_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_26_clk_i (.X(clknet_leaf_26_clk_i),
    .A(clknet_5_8__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _4886_ (.A(raddr_a_i[1]),
    .B_N(raddr_a_i[2]),
    .Y(_1002_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_25_clk_i (.X(clknet_leaf_25_clk_i),
    .A(clknet_5_8__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_24_clk_i (.X(clknet_leaf_24_clk_i),
    .A(clknet_5_8__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_23_clk_i (.X(clknet_leaf_23_clk_i),
    .A(clknet_5_9__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_22_clk_i (.X(clknet_leaf_22_clk_i),
    .A(clknet_5_9__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4891_ (.A0(rf_reg[415]),
    .A1(rf_reg[447]),
    .S(raddr_a_i[0]),
    .X(_1007_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4892_ (.Y(_1008_),
    .B1(net261),
    .B2(_1007_),
    .A2(_1000_),
    .A1(net277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4893_ (.A0(rf_reg[287]),
    .A1(rf_reg[319]),
    .S(raddr_a_i[0]),
    .X(_1009_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _4894_ (.A(raddr_a_i[1]),
    .B(raddr_a_i[2]),
    .Y(_1010_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_21_clk_i (.X(clknet_leaf_21_clk_i),
    .A(clknet_5_9__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_20_clk_i (.X(clknet_leaf_20_clk_i),
    .A(clknet_5_9__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4897_ (.A0(rf_reg[351]),
    .A1(rf_reg[383]),
    .S(raddr_a_i[0]),
    .X(_1013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _4898_ (.A(raddr_a_i[2]),
    .B_N(raddr_a_i[1]),
    .Y(_1014_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_19_clk_i (.X(clknet_leaf_19_clk_i),
    .A(clknet_5_12__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_18_clk_i (.X(clknet_leaf_18_clk_i),
    .A(clknet_5_12__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4901_ (.Y(_1017_),
    .B1(_1013_),
    .B2(net239),
    .A2(net250),
    .A1(_1009_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _4902_ (.VDD(VDD),
    .Y(_1018_),
    .A(raddr_a_i[4]),
    .VSS(VSS));
 sg13g2_nand2_1 _4903_ (.Y(_1019_),
    .A(_1018_),
    .B(raddr_a_i[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_17_clk_i (.X(clknet_leaf_17_clk_i),
    .A(clknet_5_12__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 _4905_ (.A2(_1017_),
    .A1(_1008_),
    .B1(net233),
    .X(_1021_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_16_clk_i (.X(clknet_leaf_16_clk_i),
    .A(clknet_5_13__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_15_clk_i (.X(clknet_leaf_15_clk_i),
    .A(clknet_5_6__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_14_clk_i (.X(clknet_leaf_14_clk_i),
    .A(clknet_5_6__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_13_clk_i (.X(clknet_leaf_13_clk_i),
    .A(clknet_5_6__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4910_ (.A0(rf_reg[63]),
    .A1(rf_reg[127]),
    .S(raddr_a_i[1]),
    .X(_1026_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _4911_ (.Y(_1027_),
    .A(raddr_a_i[0]),
    .B(_1026_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_12_clk_i (.X(clknet_leaf_12_clk_i),
    .A(clknet_5_3__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_11_clk_i (.X(clknet_leaf_11_clk_i),
    .A(clknet_5_3__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_10_clk_i (.X(clknet_leaf_10_clk_i),
    .A(clknet_5_3__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_9_clk_i (.X(clknet_leaf_9_clk_i),
    .A(clknet_5_3__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_8_clk_i (.X(clknet_leaf_8_clk_i),
    .A(clknet_5_2__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_7_clk_i (.X(clknet_leaf_7_clk_i),
    .A(clknet_5_2__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _4918_ (.B(rf_reg[95]),
    .C(raddr_a_i[1]),
    .Y(_1034_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_buf_16 clkbuf_leaf_6_clk_i (.X(clknet_leaf_6_clk_i),
    .A(clknet_5_2__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _4920_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1027_),
    .A2(_1034_),
    .Y(_1036_),
    .B1(raddr_a_i[2]));
 sg13g2_buf_16 clkbuf_leaf_5_clk_i (.X(clknet_leaf_5_clk_i),
    .A(clknet_5_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_4_clk_i (.X(clknet_leaf_4_clk_i),
    .A(clknet_5_2__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4923_ (.A0(rf_reg[159]),
    .A1(rf_reg[191]),
    .S(raddr_a_i[0]),
    .X(_1039_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_3_clk_i (.X(clknet_leaf_3_clk_i),
    .A(clknet_5_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4925_ (.A0(rf_reg[223]),
    .A1(rf_reg[255]),
    .S(raddr_a_i[0]),
    .X(_1041_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4926_ (.Y(_1042_),
    .B1(_1041_),
    .B2(net281),
    .A2(_1039_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _4927_ (.VDD(VDD),
    .Y(_1043_),
    .A(_1042_),
    .VSS(VSS));
 sg13g2_nor2_1 _4928_ (.A(raddr_a_i[4]),
    .B(raddr_a_i[3]),
    .Y(_1044_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_2_clk_i (.X(clknet_leaf_2_clk_i),
    .A(clknet_5_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _4930_ (.B1(net312),
    .VDD(VDD),
    .Y(_1046_),
    .VSS(VSS),
    .A1(_1036_),
    .A2(_1043_));
 sg13g2_inv_1 _4931_ (.VDD(VDD),
    .Y(_1047_),
    .A(raddr_a_i[2]),
    .VSS(VSS));
 sg13g2_nor3_1 _4932_ (.A(_1018_),
    .B(raddr_a_i[3]),
    .C(_1047_),
    .Y(_1048_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_1_clk_i (.X(clknet_leaf_1_clk_i),
    .A(clknet_5_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_0_clk_i (.X(clknet_leaf_0_clk_i),
    .A(clknet_5_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _4935_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[671]),
    .A1(rf_reg[703]),
    .A2(rf_reg[735]),
    .A3(rf_reg[767]),
    .S1(raddr_a_i[1]),
    .X(_1051_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _4936_ (.A(_1018_),
    .B(raddr_a_i[3]),
    .C(raddr_a_i[2]),
    .Y(_1052_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout315 (.A(_1044_),
    .X(net315),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _4938_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[543]),
    .A1(rf_reg[575]),
    .A2(rf_reg[607]),
    .A3(rf_reg[639]),
    .S1(raddr_a_i[1]),
    .X(_1054_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net315),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net314),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4941_ (.A0(rf_reg[991]),
    .A1(rf_reg[1023]),
    .S(raddr_a_i[0]),
    .X(_1057_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(net315),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4943_ (.A0(rf_reg[927]),
    .A1(rf_reg[959]),
    .S(raddr_a_i[0]),
    .X(_1059_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(net312),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4945_ (.Y(_1061_),
    .B1(_1059_),
    .B2(net262),
    .A2(_1057_),
    .A1(net278),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout310 (.A(_1068_),
    .X(net310),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net310),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4948_ (.A0(rf_reg[863]),
    .A1(rf_reg[895]),
    .S(raddr_a_i[0]),
    .X(_1064_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4950_ (.A0(rf_reg[799]),
    .A1(rf_reg[831]),
    .S(raddr_a_i[0]),
    .X(_1066_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4951_ (.Y(_1067_),
    .B1(_1066_),
    .B2(net250),
    .A2(_1064_),
    .A1(net239),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _4952_ (.Y(_1068_),
    .A(raddr_a_i[4]),
    .B(raddr_a_i[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _4953_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net307),
    .Y(_1069_),
    .A2(_1067_),
    .A1(_1061_));
 sg13g2_a221oi_1 _4954_ (.VSS(VSS),
    .VDD(VDD),
    .B2(_1054_),
    .C1(_1069_),
    .B1(net228),
    .A1(net67),
    .Y(_1070_),
    .A2(_1051_));
 sg13g2_nand3_1 _4955_ (.B(_1046_),
    .C(_1070_),
    .A(_1021_),
    .Y(rdata_a_o[31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4956_ (.A0(rf_reg[926]),
    .A1(rf_reg[958]),
    .S(raddr_a_i[0]),
    .X(_1071_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(net310),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4958_ (.A0(rf_reg[990]),
    .A1(rf_reg[1022]),
    .S(raddr_a_i[0]),
    .X(_1073_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(net307),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4960_ (.Y(_1075_),
    .B1(_1073_),
    .B2(net278),
    .A2(_1071_),
    .A1(net262),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(_1971_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4962_ (.A0(rf_reg[798]),
    .A1(rf_reg[830]),
    .S(raddr_a_i[0]),
    .X(_1077_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4963_ (.A0(rf_reg[862]),
    .A1(rf_reg[894]),
    .S(raddr_a_i[0]),
    .X(_1078_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4964_ (.Y(_1079_),
    .B1(_1078_),
    .B2(net240),
    .A2(_1077_),
    .A1(net251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(net305),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _4966_ (.A2(_1079_),
    .A1(_1075_),
    .B1(net307),
    .X(_1081_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4967_ (.A0(rf_reg[62]),
    .A1(rf_reg[126]),
    .S(raddr_a_i[1]),
    .X(_1082_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _4968_ (.Y(_1083_),
    .A(raddr_a_i[0]),
    .B(_1082_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _4969_ (.B(rf_reg[94]),
    .C(raddr_a_i[1]),
    .Y(_1084_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _4970_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1083_),
    .A2(_1084_),
    .Y(_1085_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _4971_ (.A0(rf_reg[158]),
    .A1(rf_reg[190]),
    .S(raddr_a_i[0]),
    .X(_1086_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(net304),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4973_ (.A0(rf_reg[222]),
    .A1(rf_reg[254]),
    .S(raddr_a_i[0]),
    .X(_1088_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4974_ (.Y(_1089_),
    .B1(_1088_),
    .B2(net281),
    .A2(_1086_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _4975_ (.VDD(VDD),
    .Y(_1090_),
    .A(_1089_),
    .VSS(VSS));
 sg13g2_o21ai_1 _4976_ (.B1(net312),
    .VDD(VDD),
    .Y(_1091_),
    .VSS(VSS),
    .A1(_1085_),
    .A2(_1090_));
 sg13g2_mux4_1 _4977_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[670]),
    .A1(rf_reg[702]),
    .A2(rf_reg[734]),
    .A3(rf_reg[766]),
    .S1(raddr_a_i[1]),
    .X(_1092_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(net305),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _4980_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[542]),
    .A1(rf_reg[574]),
    .A2(rf_reg[606]),
    .A3(rf_reg[638]),
    .S1(raddr_a_i[1]),
    .X(_1095_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4981_ (.A0(rf_reg[478]),
    .A1(rf_reg[510]),
    .S(raddr_a_i[0]),
    .X(_1096_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4982_ (.A0(rf_reg[414]),
    .A1(rf_reg[446]),
    .S(raddr_a_i[0]),
    .X(_1097_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4983_ (.Y(_1098_),
    .B1(_1097_),
    .B2(net262),
    .A2(_1096_),
    .A1(net278),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4984_ (.A0(rf_reg[350]),
    .A1(rf_reg[382]),
    .S(raddr_a_i[0]),
    .X(_1099_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4985_ (.A0(rf_reg[286]),
    .A1(rf_reg[318]),
    .S(raddr_a_i[0]),
    .X(_1100_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4986_ (.Y(_1101_),
    .B1(_1100_),
    .B2(net251),
    .A2(_1099_),
    .A1(net240),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _4987_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1098_),
    .A2(_1101_),
    .Y(_1102_),
    .B1(net233));
 sg13g2_a221oi_1 _4988_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net228),
    .C1(_1102_),
    .B1(_1095_),
    .A1(net67),
    .Y(_1103_),
    .A2(_1092_));
 sg13g2_nand3_1 _4989_ (.B(_1091_),
    .C(_1103_),
    .A(_1081_),
    .Y(rdata_a_o[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4990_ (.A0(rf_reg[917]),
    .A1(rf_reg[949]),
    .S(raddr_a_i[0]),
    .X(_1104_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout300 (.A(_2019_),
    .X(net300),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4992_ (.A0(rf_reg[981]),
    .A1(rf_reg[1013]),
    .S(raddr_a_i[0]),
    .X(_1106_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4993_ (.Y(_1107_),
    .B1(_1106_),
    .B2(net276),
    .A2(_1104_),
    .A1(net260),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4994_ (.A0(rf_reg[789]),
    .A1(rf_reg[821]),
    .S(raddr_a_i[0]),
    .X(_1108_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4995_ (.A0(rf_reg[853]),
    .A1(rf_reg[885]),
    .S(raddr_a_i[0]),
    .X(_1109_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _4996_ (.Y(_1110_),
    .B1(_1109_),
    .B2(net237),
    .A2(_1108_),
    .A1(net248),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _4997_ (.A2(_1110_),
    .A1(_1107_),
    .B1(net307),
    .X(_1111_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _4998_ (.A0(rf_reg[53]),
    .A1(rf_reg[117]),
    .S(raddr_a_i[1]),
    .X(_1112_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _4999_ (.Y(_1113_),
    .A(raddr_a_i[0]),
    .B(_1112_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5000_ (.B(rf_reg[85]),
    .C(raddr_a_i[1]),
    .Y(_1114_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5001_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1113_),
    .A2(_1114_),
    .Y(_1115_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5002_ (.A0(rf_reg[149]),
    .A1(rf_reg[181]),
    .S(raddr_a_i[0]),
    .X(_1116_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5003_ (.A0(rf_reg[213]),
    .A1(rf_reg[245]),
    .S(raddr_a_i[0]),
    .X(_1117_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5004_ (.Y(_1118_),
    .B1(_1117_),
    .B2(net280),
    .A2(_1116_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5005_ (.VDD(VDD),
    .Y(_1119_),
    .A(_1118_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5006_ (.B1(net311),
    .VDD(VDD),
    .Y(_1120_),
    .VSS(VSS),
    .A1(_1115_),
    .A2(_1119_));
 sg13g2_mux4_1 _5007_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[661]),
    .A1(rf_reg[693]),
    .A2(rf_reg[725]),
    .A3(rf_reg[757]),
    .S1(raddr_a_i[1]),
    .X(_1121_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5008_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[533]),
    .A1(rf_reg[565]),
    .A2(rf_reg[597]),
    .A3(rf_reg[629]),
    .S1(raddr_a_i[1]),
    .X(_1122_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5009_ (.A0(rf_reg[469]),
    .A1(rf_reg[501]),
    .S(raddr_a_i[0]),
    .X(_1123_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5010_ (.A0(rf_reg[405]),
    .A1(rf_reg[437]),
    .S(raddr_a_i[0]),
    .X(_1124_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5011_ (.Y(_1125_),
    .B1(_1124_),
    .B2(net260),
    .A2(_1123_),
    .A1(net276),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5012_ (.A0(rf_reg[341]),
    .A1(rf_reg[373]),
    .S(raddr_a_i[0]),
    .X(_1126_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5013_ (.A0(rf_reg[277]),
    .A1(rf_reg[309]),
    .S(raddr_a_i[0]),
    .X(_1127_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5014_ (.Y(_1128_),
    .B1(_1127_),
    .B2(net248),
    .A2(_1126_),
    .A1(net237),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5015_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1125_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(net232));
 sg13g2_a221oi_1 _5016_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1129_),
    .B1(_1122_),
    .A1(net66),
    .Y(_1130_),
    .A2(_1121_));
 sg13g2_nand3_1 _5017_ (.B(_1120_),
    .C(_1130_),
    .A(_1111_),
    .Y(rdata_a_o[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5018_ (.A0(rf_reg[916]),
    .A1(rf_reg[948]),
    .S(raddr_a_i[0]),
    .X(_1131_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5019_ (.A0(rf_reg[980]),
    .A1(rf_reg[1012]),
    .S(raddr_a_i[0]),
    .X(_1132_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5020_ (.Y(_1133_),
    .B1(_1132_),
    .B2(net285),
    .A2(_1131_),
    .A1(net269),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(net300),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5022_ (.A0(rf_reg[788]),
    .A1(rf_reg[820]),
    .S(raddr_a_i[0]),
    .X(_1135_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5023_ (.A0(rf_reg[852]),
    .A1(rf_reg[884]),
    .S(raddr_a_i[0]),
    .X(_1136_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5024_ (.Y(_1137_),
    .B1(_1136_),
    .B2(net244),
    .A2(_1135_),
    .A1(net255),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5025_ (.A2(_1137_),
    .A1(_1133_),
    .B1(net308),
    .X(_1138_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5026_ (.A0(rf_reg[52]),
    .A1(rf_reg[116]),
    .S(raddr_a_i[1]),
    .X(_1139_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5027_ (.Y(_1140_),
    .A(raddr_a_i[0]),
    .B(_1139_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5028_ (.B(rf_reg[84]),
    .C(raddr_a_i[1]),
    .Y(_1141_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5029_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1140_),
    .A2(_1141_),
    .Y(_1142_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5030_ (.A0(rf_reg[148]),
    .A1(rf_reg[180]),
    .S(raddr_a_i[0]),
    .X(_1143_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5031_ (.A0(rf_reg[212]),
    .A1(rf_reg[244]),
    .S(raddr_a_i[0]),
    .X(_1144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5032_ (.Y(_1145_),
    .B1(_1144_),
    .B2(net288),
    .A2(_1143_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5033_ (.VDD(VDD),
    .Y(_1146_),
    .A(_1145_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5034_ (.B1(net313),
    .VDD(VDD),
    .Y(_1147_),
    .VSS(VSS),
    .A1(_1142_),
    .A2(_1146_));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5036_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[660]),
    .A1(rf_reg[692]),
    .A2(rf_reg[724]),
    .A3(rf_reg[756]),
    .S1(raddr_a_i[1]),
    .X(_1149_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5037_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[532]),
    .A1(rf_reg[564]),
    .A2(rf_reg[596]),
    .A3(rf_reg[628]),
    .S1(raddr_a_i[1]),
    .X(_1150_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5038_ (.A0(rf_reg[468]),
    .A1(rf_reg[500]),
    .S(raddr_a_i[0]),
    .X(_1151_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5039_ (.A0(rf_reg[404]),
    .A1(rf_reg[436]),
    .S(raddr_a_i[0]),
    .X(_1152_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5040_ (.Y(_1153_),
    .B1(_1152_),
    .B2(net269),
    .A2(_1151_),
    .A1(net285),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5041_ (.A0(rf_reg[340]),
    .A1(rf_reg[372]),
    .S(raddr_a_i[0]),
    .X(_1154_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5042_ (.A0(rf_reg[276]),
    .A1(rf_reg[308]),
    .S(raddr_a_i[0]),
    .X(_1155_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5043_ (.Y(_1156_),
    .B1(_1155_),
    .B2(net255),
    .A2(_1154_),
    .A1(net244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5044_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net234),
    .Y(_1157_),
    .A2(_1156_),
    .A1(_1153_));
 sg13g2_a221oi_1 _5045_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1157_),
    .B1(_1150_),
    .A1(net68),
    .Y(_1158_),
    .A2(_1149_));
 sg13g2_nand3_1 _5046_ (.B(_1147_),
    .C(_1158_),
    .A(_1138_),
    .Y(rdata_a_o[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5047_ (.A0(rf_reg[915]),
    .A1(rf_reg[947]),
    .S(raddr_a_i[0]),
    .X(_1159_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5048_ (.A0(rf_reg[979]),
    .A1(rf_reg[1011]),
    .S(raddr_a_i[0]),
    .X(_1160_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5049_ (.Y(_1161_),
    .B1(_1160_),
    .B2(net284),
    .A2(_1159_),
    .A1(net268),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5050_ (.A0(rf_reg[787]),
    .A1(rf_reg[819]),
    .S(raddr_a_i[0]),
    .X(_1162_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5051_ (.A0(rf_reg[851]),
    .A1(rf_reg[883]),
    .S(raddr_a_i[0]),
    .X(_1163_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5052_ (.Y(_1164_),
    .B1(_1163_),
    .B2(net243),
    .A2(_1162_),
    .A1(net254),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5053_ (.A2(_1164_),
    .A1(_1161_),
    .B1(net309),
    .X(_1165_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5054_ (.A0(rf_reg[51]),
    .A1(rf_reg[115]),
    .S(raddr_a_i[1]),
    .X(_1166_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5055_ (.Y(_1167_),
    .A(raddr_a_i[0]),
    .B(_1166_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5056_ (.B(rf_reg[83]),
    .C(raddr_a_i[1]),
    .Y(_1168_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5057_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1167_),
    .A2(_1168_),
    .Y(_1169_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5058_ (.A0(rf_reg[147]),
    .A1(rf_reg[179]),
    .S(raddr_a_i[0]),
    .X(_1170_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5059_ (.A0(rf_reg[211]),
    .A1(rf_reg[243]),
    .S(raddr_a_i[0]),
    .X(_1171_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5060_ (.Y(_1172_),
    .B1(_1171_),
    .B2(net289),
    .A2(_1170_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5061_ (.VDD(VDD),
    .Y(_1173_),
    .A(_1172_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5062_ (.B1(net314),
    .VDD(VDD),
    .Y(_1174_),
    .VSS(VSS),
    .A1(_1169_),
    .A2(_1173_));
 sg13g2_mux4_1 _5063_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[659]),
    .A1(rf_reg[691]),
    .A2(rf_reg[723]),
    .A3(rf_reg[755]),
    .S1(raddr_a_i[1]),
    .X(_1175_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5064_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[531]),
    .A1(rf_reg[563]),
    .A2(rf_reg[595]),
    .A3(rf_reg[627]),
    .S1(raddr_a_i[1]),
    .X(_1176_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5065_ (.A0(rf_reg[467]),
    .A1(rf_reg[499]),
    .S(raddr_a_i[0]),
    .X(_1177_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5066_ (.A0(rf_reg[403]),
    .A1(rf_reg[435]),
    .S(raddr_a_i[0]),
    .X(_1178_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5067_ (.Y(_1179_),
    .B1(_1178_),
    .B2(net268),
    .A2(_1177_),
    .A1(net284),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5068_ (.A0(rf_reg[339]),
    .A1(rf_reg[371]),
    .S(raddr_a_i[0]),
    .X(_1180_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5069_ (.A0(rf_reg[275]),
    .A1(rf_reg[307]),
    .S(raddr_a_i[0]),
    .X(_1181_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5070_ (.Y(_1182_),
    .B1(_1181_),
    .B2(net254),
    .A2(_1180_),
    .A1(net243),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5071_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1179_),
    .A2(_1182_),
    .Y(_1183_),
    .B1(net235));
 sg13g2_a221oi_1 _5072_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1183_),
    .B1(_1176_),
    .A1(net69),
    .Y(_1184_),
    .A2(_1175_));
 sg13g2_nand3_1 _5073_ (.B(_1174_),
    .C(_1184_),
    .A(_1165_),
    .Y(rdata_a_o[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5074_ (.A0(rf_reg[914]),
    .A1(rf_reg[946]),
    .S(raddr_a_i[0]),
    .X(_1185_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5075_ (.A0(rf_reg[978]),
    .A1(rf_reg[1010]),
    .S(raddr_a_i[0]),
    .X(_1186_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5076_ (.Y(_1187_),
    .B1(_1186_),
    .B2(net284),
    .A2(_1185_),
    .A1(net267),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5077_ (.A0(rf_reg[786]),
    .A1(rf_reg[818]),
    .S(raddr_a_i[0]),
    .X(_1188_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5078_ (.A0(rf_reg[850]),
    .A1(rf_reg[882]),
    .S(raddr_a_i[0]),
    .X(_1189_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5079_ (.Y(_1190_),
    .B1(_1189_),
    .B2(net242),
    .A2(_1188_),
    .A1(net254),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5080_ (.A2(_1190_),
    .A1(_1187_),
    .B1(net309),
    .X(_1191_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net300),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5082_ (.A0(rf_reg[50]),
    .A1(rf_reg[114]),
    .S(raddr_a_i[1]),
    .X(_1193_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5083_ (.Y(_1194_),
    .A(raddr_a_i[0]),
    .B(_1193_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5084_ (.B(rf_reg[82]),
    .C(raddr_a_i[1]),
    .Y(_1195_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5085_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1194_),
    .A2(_1195_),
    .Y(_1196_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5086_ (.A0(rf_reg[146]),
    .A1(rf_reg[178]),
    .S(raddr_a_i[0]),
    .X(_1197_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5087_ (.A0(rf_reg[210]),
    .A1(rf_reg[242]),
    .S(raddr_a_i[0]),
    .X(_1198_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5088_ (.Y(_1199_),
    .B1(_1198_),
    .B2(net289),
    .A2(_1197_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5089_ (.VDD(VDD),
    .Y(_1200_),
    .A(_1199_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5090_ (.B1(net314),
    .VDD(VDD),
    .Y(_1201_),
    .VSS(VSS),
    .A1(_1196_),
    .A2(_1200_));
 sg13g2_mux4_1 _5091_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[658]),
    .A1(rf_reg[690]),
    .A2(rf_reg[722]),
    .A3(rf_reg[754]),
    .S1(raddr_a_i[1]),
    .X(_1202_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5092_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[530]),
    .A1(rf_reg[562]),
    .A2(rf_reg[594]),
    .A3(rf_reg[626]),
    .S1(raddr_a_i[1]),
    .X(_1203_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5093_ (.A0(rf_reg[466]),
    .A1(rf_reg[498]),
    .S(raddr_a_i[0]),
    .X(_1204_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5094_ (.A0(rf_reg[402]),
    .A1(rf_reg[434]),
    .S(raddr_a_i[0]),
    .X(_1205_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5095_ (.Y(_1206_),
    .B1(_1205_),
    .B2(net268),
    .A2(_1204_),
    .A1(net284),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5096_ (.A0(rf_reg[338]),
    .A1(rf_reg[370]),
    .S(raddr_a_i[0]),
    .X(_1207_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5098_ (.A0(rf_reg[274]),
    .A1(rf_reg[306]),
    .S(raddr_a_i[0]),
    .X(_1209_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5099_ (.Y(_1210_),
    .B1(_1209_),
    .B2(net254),
    .A2(_1207_),
    .A1(net243),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5100_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net235),
    .Y(_1211_),
    .A2(_1210_),
    .A1(_1206_));
 sg13g2_a221oi_1 _5101_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1211_),
    .B1(_1203_),
    .A1(net69),
    .Y(_1212_),
    .A2(_1202_));
 sg13g2_nand3_1 _5102_ (.B(_1201_),
    .C(_1212_),
    .A(_1191_),
    .Y(rdata_a_o[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5103_ (.A0(rf_reg[913]),
    .A1(rf_reg[945]),
    .S(raddr_a_i[0]),
    .X(_1213_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5104_ (.A0(rf_reg[977]),
    .A1(rf_reg[1009]),
    .S(raddr_a_i[0]),
    .X(_1214_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5105_ (.Y(_1215_),
    .B1(_1214_),
    .B2(net276),
    .A2(_1213_),
    .A1(net260),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5106_ (.A0(rf_reg[785]),
    .A1(rf_reg[817]),
    .S(raddr_a_i[0]),
    .X(_1216_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5107_ (.A0(rf_reg[849]),
    .A1(rf_reg[881]),
    .S(raddr_a_i[0]),
    .X(_1217_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5108_ (.Y(_1218_),
    .B1(_1217_),
    .B2(net237),
    .A2(_1216_),
    .A1(net248),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5109_ (.A2(_1218_),
    .A1(_1215_),
    .B1(net306),
    .X(_1219_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5110_ (.A0(rf_reg[49]),
    .A1(rf_reg[113]),
    .S(raddr_a_i[1]),
    .X(_1220_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5111_ (.Y(_1221_),
    .A(raddr_a_i[0]),
    .B(_1220_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout295 (.A(_2034_),
    .X(net295),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5113_ (.B(rf_reg[81]),
    .C(raddr_a_i[1]),
    .Y(_1223_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5114_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1221_),
    .A2(_1223_),
    .Y(_1224_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5115_ (.A0(rf_reg[145]),
    .A1(rf_reg[177]),
    .S(raddr_a_i[0]),
    .X(_1225_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5116_ (.A0(rf_reg[209]),
    .A1(rf_reg[241]),
    .S(raddr_a_i[0]),
    .X(_1226_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5117_ (.Y(_1227_),
    .B1(_1226_),
    .B2(net280),
    .A2(_1225_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5118_ (.VDD(VDD),
    .Y(_1228_),
    .A(_1227_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5119_ (.B1(net311),
    .VDD(VDD),
    .Y(_1229_),
    .VSS(VSS),
    .A1(_1224_),
    .A2(_1228_));
 sg13g2_mux4_1 _5120_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[657]),
    .A1(rf_reg[689]),
    .A2(rf_reg[721]),
    .A3(rf_reg[753]),
    .S1(raddr_a_i[1]),
    .X(_1230_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5121_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[529]),
    .A1(rf_reg[561]),
    .A2(rf_reg[593]),
    .A3(rf_reg[625]),
    .S1(raddr_a_i[1]),
    .X(_1231_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(net295),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5123_ (.A0(rf_reg[465]),
    .A1(rf_reg[497]),
    .S(raddr_a_i[0]),
    .X(_1233_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5124_ (.A0(rf_reg[401]),
    .A1(rf_reg[433]),
    .S(raddr_a_i[0]),
    .X(_1234_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net294),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5126_ (.Y(_1236_),
    .B1(_1234_),
    .B2(net260),
    .A2(_1233_),
    .A1(net276),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5127_ (.A0(rf_reg[337]),
    .A1(rf_reg[369]),
    .S(raddr_a_i[0]),
    .X(_1237_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5128_ (.A0(rf_reg[273]),
    .A1(rf_reg[305]),
    .S(raddr_a_i[0]),
    .X(_1238_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5129_ (.Y(_1239_),
    .B1(_1238_),
    .B2(net248),
    .A2(_1237_),
    .A1(net237),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5130_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net232),
    .Y(_1240_),
    .A2(_1239_),
    .A1(_1236_));
 sg13g2_a221oi_1 _5131_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1240_),
    .B1(_1231_),
    .A1(net66),
    .Y(_1241_),
    .A2(_1230_));
 sg13g2_nand3_1 _5132_ (.B(_1229_),
    .C(_1241_),
    .A(_1219_),
    .Y(rdata_a_o[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(net295),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5134_ (.A0(rf_reg[912]),
    .A1(rf_reg[944]),
    .S(raddr_a_i[0]),
    .X(_1243_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5135_ (.A0(rf_reg[976]),
    .A1(rf_reg[1008]),
    .S(raddr_a_i[0]),
    .X(_1244_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5136_ (.Y(_1245_),
    .B1(_1244_),
    .B2(net283),
    .A2(_1243_),
    .A1(net267),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5137_ (.A0(rf_reg[784]),
    .A1(rf_reg[816]),
    .S(raddr_a_i[0]),
    .X(_1246_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5138_ (.A0(rf_reg[848]),
    .A1(rf_reg[880]),
    .S(raddr_a_i[0]),
    .X(_1247_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5139_ (.Y(_1248_),
    .B1(_1247_),
    .B2(net244),
    .A2(_1246_),
    .A1(net253),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 _5140_ (.A2(_1248_),
    .A1(_1245_),
    .B1(net308),
    .X(_1249_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5141_ (.A0(rf_reg[48]),
    .A1(rf_reg[112]),
    .S(raddr_a_i[1]),
    .X(_1250_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5142_ (.Y(_1251_),
    .A(raddr_a_i[0]),
    .B(_1250_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5143_ (.B(rf_reg[80]),
    .C(raddr_a_i[1]),
    .Y(_1252_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5144_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1251_),
    .A2(_1252_),
    .Y(_1253_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5145_ (.A0(rf_reg[144]),
    .A1(rf_reg[176]),
    .S(raddr_a_i[0]),
    .X(_1254_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5146_ (.A0(rf_reg[208]),
    .A1(rf_reg[240]),
    .S(raddr_a_i[0]),
    .X(_1255_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5147_ (.Y(_1256_),
    .B1(_1255_),
    .B2(net289),
    .A2(_1254_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5148_ (.VDD(VDD),
    .Y(_1257_),
    .A(_1256_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5149_ (.B1(net313),
    .VDD(VDD),
    .Y(_1258_),
    .VSS(VSS),
    .A1(_1253_),
    .A2(_1257_));
 sg13g2_mux4_1 _5150_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[656]),
    .A1(rf_reg[688]),
    .A2(rf_reg[720]),
    .A3(rf_reg[752]),
    .S1(raddr_a_i[1]),
    .X(_1259_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(net292),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5152_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[528]),
    .A1(rf_reg[560]),
    .A2(rf_reg[592]),
    .A3(rf_reg[624]),
    .S1(raddr_a_i[1]),
    .X(_1261_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5153_ (.A0(rf_reg[464]),
    .A1(rf_reg[496]),
    .S(raddr_a_i[0]),
    .X(_1262_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(_0993_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5155_ (.A0(rf_reg[400]),
    .A1(rf_reg[432]),
    .S(raddr_a_i[0]),
    .X(_1264_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5156_ (.Y(_1265_),
    .B1(_1264_),
    .B2(net267),
    .A2(_1262_),
    .A1(net283),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5157_ (.A0(rf_reg[336]),
    .A1(rf_reg[368]),
    .S(raddr_a_i[0]),
    .X(_1266_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5158_ (.A0(rf_reg[272]),
    .A1(rf_reg[304]),
    .S(raddr_a_i[0]),
    .X(_1267_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5159_ (.Y(_1268_),
    .B1(_1267_),
    .B2(net255),
    .A2(_1266_),
    .A1(net244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5160_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net234),
    .Y(_1269_),
    .A2(_1268_),
    .A1(_1265_));
 sg13g2_a221oi_1 _5161_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1269_),
    .B1(_1261_),
    .A1(net68),
    .Y(_1270_),
    .A2(_1259_));
 sg13g2_nand3_1 _5162_ (.B(_1258_),
    .C(_1270_),
    .A(_1249_),
    .Y(rdata_a_o[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5163_ (.A0(rf_reg[911]),
    .A1(rf_reg[943]),
    .S(raddr_a_i[0]),
    .X(_1271_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5164_ (.A0(rf_reg[975]),
    .A1(rf_reg[1007]),
    .S(raddr_a_i[0]),
    .X(_1272_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5165_ (.Y(_1273_),
    .B1(_1272_),
    .B2(net278),
    .A2(_1271_),
    .A1(net262),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5166_ (.A0(rf_reg[783]),
    .A1(rf_reg[815]),
    .S(raddr_a_i[0]),
    .X(_1274_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5167_ (.A0(rf_reg[847]),
    .A1(rf_reg[879]),
    .S(raddr_a_i[0]),
    .X(_1275_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5168_ (.Y(_1276_),
    .B1(_1275_),
    .B2(net240),
    .A2(_1274_),
    .A1(net251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5169_ (.A2(_1276_),
    .A1(_1273_),
    .B1(net307),
    .X(_1277_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5170_ (.A0(rf_reg[47]),
    .A1(rf_reg[111]),
    .S(raddr_a_i[1]),
    .X(_1278_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5171_ (.Y(_1279_),
    .A(raddr_a_i[0]),
    .B(_1278_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(net290),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5173_ (.B(rf_reg[79]),
    .C(raddr_a_i[1]),
    .Y(_1281_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5174_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1279_),
    .A2(_1281_),
    .Y(_1282_),
    .B1(raddr_a_i[2]));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(net289),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5176_ (.A0(rf_reg[143]),
    .A1(rf_reg[175]),
    .S(raddr_a_i[0]),
    .X(_1284_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5177_ (.A0(rf_reg[207]),
    .A1(rf_reg[239]),
    .S(raddr_a_i[0]),
    .X(_1285_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout287 (.A(net290),
    .X(net287),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5179_ (.Y(_1287_),
    .B1(_1285_),
    .B2(net282),
    .A2(_1284_),
    .A1(net266),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5180_ (.VDD(VDD),
    .Y(_1288_),
    .A(_1287_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5181_ (.B1(net312),
    .VDD(VDD),
    .Y(_1289_),
    .VSS(VSS),
    .A1(_1282_),
    .A2(_1288_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(net287),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5183_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[655]),
    .A1(rf_reg[687]),
    .A2(rf_reg[719]),
    .A3(rf_reg[751]),
    .S1(raddr_a_i[1]),
    .X(_1291_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5184_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[527]),
    .A1(rf_reg[559]),
    .A2(rf_reg[591]),
    .A3(rf_reg[623]),
    .S1(raddr_a_i[1]),
    .X(_1292_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5185_ (.A0(rf_reg[463]),
    .A1(rf_reg[495]),
    .S(raddr_a_i[0]),
    .X(_1293_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5186_ (.A0(rf_reg[399]),
    .A1(rf_reg[431]),
    .S(raddr_a_i[0]),
    .X(_1294_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5187_ (.Y(_1295_),
    .B1(_1294_),
    .B2(net268),
    .A2(_1293_),
    .A1(net284),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net286),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net287),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5190_ (.A0(rf_reg[335]),
    .A1(rf_reg[367]),
    .S(raddr_a_i[0]),
    .X(_1298_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5191_ (.A0(rf_reg[271]),
    .A1(rf_reg[303]),
    .S(raddr_a_i[0]),
    .X(_1299_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(net287),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5193_ (.Y(_1301_),
    .B1(_1299_),
    .B2(net254),
    .A2(_1298_),
    .A1(net243),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5194_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1295_),
    .A2(_1301_),
    .Y(_1302_),
    .B1(net235));
 sg13g2_a221oi_1 _5195_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net228),
    .C1(_1302_),
    .B1(_1292_),
    .A1(net67),
    .Y(_1303_),
    .A2(_1291_));
 sg13g2_nand3_1 _5196_ (.B(_1289_),
    .C(_1303_),
    .A(_1277_),
    .Y(rdata_a_o[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5197_ (.A0(rf_reg[910]),
    .A1(rf_reg[942]),
    .S(raddr_a_i[0]),
    .X(_1304_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5198_ (.A0(rf_reg[974]),
    .A1(rf_reg[1006]),
    .S(raddr_a_i[0]),
    .X(_1305_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5199_ (.Y(_1306_),
    .B1(_1305_),
    .B2(net283),
    .A2(_1304_),
    .A1(net261),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5200_ (.A0(rf_reg[782]),
    .A1(rf_reg[814]),
    .S(raddr_a_i[0]),
    .X(_1307_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5201_ (.A0(rf_reg[846]),
    .A1(rf_reg[878]),
    .S(raddr_a_i[0]),
    .X(_1308_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5202_ (.Y(_1309_),
    .B1(_1308_),
    .B2(net242),
    .A2(_1307_),
    .A1(net253),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5203_ (.A2(_1309_),
    .A1(_1306_),
    .B1(net309),
    .X(_1310_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5204_ (.A0(rf_reg[46]),
    .A1(rf_reg[110]),
    .S(raddr_a_i[1]),
    .X(_1311_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5205_ (.Y(_1312_),
    .A(raddr_a_i[0]),
    .B(_1311_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5206_ (.B(rf_reg[78]),
    .C(raddr_a_i[1]),
    .Y(_1313_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5207_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1312_),
    .A2(_1313_),
    .Y(_1314_),
    .B1(raddr_a_i[2]));
 sg13g2_buf_2 fanout282 (.A(net290),
    .X(net282),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5209_ (.A0(rf_reg[142]),
    .A1(rf_reg[174]),
    .S(raddr_a_i[0]),
    .X(_1316_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5210_ (.A0(rf_reg[206]),
    .A1(rf_reg[238]),
    .S(raddr_a_i[0]),
    .X(_1317_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5211_ (.Y(_1318_),
    .B1(_1317_),
    .B2(net281),
    .A2(_1316_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5212_ (.VDD(VDD),
    .Y(_1319_),
    .A(_1318_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5213_ (.B1(net312),
    .VDD(VDD),
    .Y(_1320_),
    .VSS(VSS),
    .A1(_1314_),
    .A2(_1319_));
 sg13g2_mux4_1 _5214_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[654]),
    .A1(rf_reg[686]),
    .A2(rf_reg[718]),
    .A3(rf_reg[750]),
    .S1(raddr_a_i[1]),
    .X(_1321_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5215_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[526]),
    .A1(rf_reg[558]),
    .A2(rf_reg[590]),
    .A3(rf_reg[622]),
    .S1(raddr_a_i[1]),
    .X(_1322_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5216_ (.A0(rf_reg[462]),
    .A1(rf_reg[494]),
    .S(raddr_a_i[0]),
    .X(_1323_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5217_ (.A0(rf_reg[398]),
    .A1(rf_reg[430]),
    .S(raddr_a_i[0]),
    .X(_1324_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5218_ (.Y(_1325_),
    .B1(_1324_),
    .B2(net262),
    .A2(_1323_),
    .A1(net277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5219_ (.A0(rf_reg[334]),
    .A1(rf_reg[366]),
    .S(raddr_a_i[0]),
    .X(_1326_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5220_ (.A0(rf_reg[270]),
    .A1(rf_reg[302]),
    .S(raddr_a_i[0]),
    .X(_1327_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5221_ (.Y(_1328_),
    .B1(_1327_),
    .B2(net251),
    .A2(_1326_),
    .A1(net240),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5222_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net233),
    .Y(_1329_),
    .A2(_1328_),
    .A1(_1325_));
 sg13g2_a221oi_1 _5223_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net228),
    .C1(_1329_),
    .B1(_1322_),
    .A1(net67),
    .Y(_1330_),
    .A2(_1321_));
 sg13g2_nand3_1 _5224_ (.B(_1320_),
    .C(_1330_),
    .A(_1310_),
    .Y(rdata_a_o[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net282),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5226_ (.A0(rf_reg[909]),
    .A1(rf_reg[941]),
    .S(raddr_a_i[0]),
    .X(_1332_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5227_ (.A0(rf_reg[973]),
    .A1(rf_reg[1005]),
    .S(raddr_a_i[0]),
    .X(_1333_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5228_ (.Y(_1334_),
    .B1(_1333_),
    .B2(net285),
    .A2(_1332_),
    .A1(net269),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5229_ (.A0(rf_reg[781]),
    .A1(rf_reg[813]),
    .S(raddr_a_i[0]),
    .X(_1335_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net281),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5231_ (.A0(rf_reg[845]),
    .A1(rf_reg[877]),
    .S(raddr_a_i[0]),
    .X(_1337_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout279 (.A(net282),
    .X(net279),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5233_ (.Y(_1339_),
    .B1(_1337_),
    .B2(net244),
    .A2(_1335_),
    .A1(net255),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5234_ (.A2(_1339_),
    .A1(_1334_),
    .B1(net308),
    .X(_1340_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net279),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5236_ (.A0(rf_reg[45]),
    .A1(rf_reg[109]),
    .S(raddr_a_i[1]),
    .X(_1342_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5237_ (.Y(_1343_),
    .A(raddr_a_i[0]),
    .B(_1342_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5238_ (.B(rf_reg[77]),
    .C(raddr_a_i[1]),
    .Y(_1344_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net279),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5240_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1343_),
    .A2(_1344_),
    .Y(_1346_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5241_ (.A0(rf_reg[141]),
    .A1(rf_reg[173]),
    .S(raddr_a_i[0]),
    .X(_1347_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5242_ (.A0(rf_reg[205]),
    .A1(rf_reg[237]),
    .S(raddr_a_i[0]),
    .X(_1348_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5243_ (.Y(_1349_),
    .B1(_1348_),
    .B2(net288),
    .A2(_1347_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5244_ (.VDD(VDD),
    .Y(_1350_),
    .A(_1349_),
    .VSS(VSS));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net279),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _5246_ (.B1(net313),
    .VDD(VDD),
    .Y(_1352_),
    .VSS(VSS),
    .A1(_1346_),
    .A2(_1350_));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(net279),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5248_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[653]),
    .A1(rf_reg[685]),
    .A2(rf_reg[717]),
    .A3(rf_reg[749]),
    .S1(raddr_a_i[1]),
    .X(_1354_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5249_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[525]),
    .A1(rf_reg[557]),
    .A2(rf_reg[589]),
    .A3(rf_reg[621]),
    .S1(raddr_a_i[1]),
    .X(_1355_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_1002_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(net274),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5252_ (.A0(rf_reg[461]),
    .A1(rf_reg[493]),
    .S(raddr_a_i[0]),
    .X(_1358_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5253_ (.A0(rf_reg[397]),
    .A1(rf_reg[429]),
    .S(raddr_a_i[0]),
    .X(_1359_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5254_ (.Y(_1360_),
    .B1(_1359_),
    .B2(net269),
    .A2(_1358_),
    .A1(net285),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5255_ (.A0(rf_reg[333]),
    .A1(rf_reg[365]),
    .S(raddr_a_i[0]),
    .X(_1361_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5256_ (.A0(rf_reg[269]),
    .A1(rf_reg[301]),
    .S(raddr_a_i[0]),
    .X(_1362_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5257_ (.Y(_1363_),
    .B1(_1362_),
    .B2(net255),
    .A2(_1361_),
    .A1(net244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5259_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net234),
    .Y(_1365_),
    .A2(_1363_),
    .A1(_1360_));
 sg13g2_a221oi_1 _5260_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1365_),
    .B1(_1355_),
    .A1(net68),
    .Y(_1366_),
    .A2(_1354_));
 sg13g2_nand3_1 _5261_ (.B(_1352_),
    .C(_1366_),
    .A(_1340_),
    .Y(rdata_a_o[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5262_ (.A0(rf_reg[908]),
    .A1(rf_reg[940]),
    .S(raddr_a_i[0]),
    .X(_1367_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5263_ (.A0(rf_reg[972]),
    .A1(rf_reg[1004]),
    .S(raddr_a_i[0]),
    .X(_1368_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout271 (.A(net274),
    .X(net271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5265_ (.Y(_1370_),
    .B1(_1368_),
    .B2(net277),
    .A2(_1367_),
    .A1(net261),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5267_ (.A0(rf_reg[780]),
    .A1(rf_reg[812]),
    .S(raddr_a_i[0]),
    .X(_1372_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5268_ (.A0(rf_reg[844]),
    .A1(rf_reg[876]),
    .S(raddr_a_i[0]),
    .X(_1373_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5269_ (.Y(_1374_),
    .B1(_1373_),
    .B2(net239),
    .A2(_1372_),
    .A1(net250),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net270),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5271_ (.A2(_1374_),
    .A1(_1370_),
    .B1(net307),
    .X(_1376_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5272_ (.A0(rf_reg[44]),
    .A1(rf_reg[108]),
    .S(raddr_a_i[1]),
    .X(_1377_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5273_ (.Y(_1378_),
    .A(raddr_a_i[0]),
    .B(_1377_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5274_ (.B(rf_reg[76]),
    .C(raddr_a_i[1]),
    .Y(_1379_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5275_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1378_),
    .A2(_1379_),
    .Y(_1380_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5276_ (.A0(rf_reg[140]),
    .A1(rf_reg[172]),
    .S(raddr_a_i[0]),
    .X(_1381_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5278_ (.A0(rf_reg[204]),
    .A1(rf_reg[236]),
    .S(raddr_a_i[0]),
    .X(_1383_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5279_ (.Y(_1384_),
    .B1(_1383_),
    .B2(net281),
    .A2(_1381_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5280_ (.VDD(VDD),
    .Y(_1385_),
    .A(_1384_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5281_ (.B1(net315),
    .VDD(VDD),
    .Y(_1386_),
    .VSS(VSS),
    .A1(_1380_),
    .A2(_1385_));
 sg13g2_mux4_1 _5282_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[652]),
    .A1(rf_reg[684]),
    .A2(rf_reg[716]),
    .A3(rf_reg[748]),
    .S1(raddr_a_i[1]),
    .X(_1387_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(net271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5284_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[524]),
    .A1(rf_reg[556]),
    .A2(rf_reg[588]),
    .A3(rf_reg[620]),
    .S1(raddr_a_i[1]),
    .X(_1389_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5285_ (.A0(rf_reg[460]),
    .A1(rf_reg[492]),
    .S(raddr_a_i[0]),
    .X(_1390_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5286_ (.A0(rf_reg[396]),
    .A1(rf_reg[428]),
    .S(raddr_a_i[0]),
    .X(_1391_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5287_ (.Y(_1392_),
    .B1(_1391_),
    .B2(net261),
    .A2(_1390_),
    .A1(net277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5288_ (.A0(rf_reg[332]),
    .A1(rf_reg[364]),
    .S(raddr_a_i[0]),
    .X(_1393_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5289_ (.A0(rf_reg[268]),
    .A1(rf_reg[300]),
    .S(raddr_a_i[0]),
    .X(_1394_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5290_ (.Y(_1395_),
    .B1(_1394_),
    .B2(net250),
    .A2(_1393_),
    .A1(net239),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5291_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net233),
    .Y(_1396_),
    .A2(_1395_),
    .A1(_1392_));
 sg13g2_a221oi_1 _5292_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net231),
    .C1(_1396_),
    .B1(_1389_),
    .A1(net70),
    .Y(_1397_),
    .A2(_1387_));
 sg13g2_nand3_1 _5293_ (.B(_1386_),
    .C(_1397_),
    .A(_1376_),
    .Y(rdata_a_o[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5294_ (.A0(rf_reg[925]),
    .A1(rf_reg[957]),
    .S(raddr_a_i[0]),
    .X(_1398_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout266 (.A(net274),
    .X(net266),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5296_ (.A0(rf_reg[989]),
    .A1(rf_reg[1021]),
    .S(raddr_a_i[0]),
    .X(_1400_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5297_ (.Y(_1401_),
    .B1(_1400_),
    .B2(net276),
    .A2(_1398_),
    .A1(net260),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5298_ (.A0(rf_reg[797]),
    .A1(rf_reg[829]),
    .S(raddr_a_i[0]),
    .X(_1402_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5299_ (.A0(rf_reg[861]),
    .A1(rf_reg[893]),
    .S(raddr_a_i[0]),
    .X(_1403_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5300_ (.Y(_1404_),
    .B1(_1403_),
    .B2(net237),
    .A2(_1402_),
    .A1(net248),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5301_ (.A2(_1404_),
    .A1(_1401_),
    .B1(net306),
    .X(_1405_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5302_ (.A0(rf_reg[61]),
    .A1(rf_reg[125]),
    .S(raddr_a_i[1]),
    .X(_1406_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5303_ (.Y(_1407_),
    .A(raddr_a_i[0]),
    .B(_1406_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5304_ (.B(rf_reg[93]),
    .C(raddr_a_i[1]),
    .Y(_1408_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5305_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1407_),
    .A2(_1408_),
    .Y(_1409_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5306_ (.A0(rf_reg[157]),
    .A1(rf_reg[189]),
    .S(raddr_a_i[0]),
    .X(_1410_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5307_ (.A0(rf_reg[221]),
    .A1(rf_reg[253]),
    .S(raddr_a_i[0]),
    .X(_1411_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5308_ (.Y(_1412_),
    .B1(_1411_),
    .B2(net280),
    .A2(_1410_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5309_ (.VDD(VDD),
    .Y(_1413_),
    .A(_1412_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5310_ (.B1(net311),
    .VDD(VDD),
    .Y(_1414_),
    .VSS(VSS),
    .A1(_1409_),
    .A2(_1413_));
 sg13g2_mux4_1 _5311_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[669]),
    .A1(rf_reg[701]),
    .A2(rf_reg[733]),
    .A3(rf_reg[765]),
    .S1(raddr_a_i[1]),
    .X(_1415_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5312_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[541]),
    .A1(rf_reg[573]),
    .A2(rf_reg[605]),
    .A3(rf_reg[637]),
    .S1(raddr_a_i[1]),
    .X(_1416_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5313_ (.A0(rf_reg[477]),
    .A1(rf_reg[509]),
    .S(raddr_a_i[0]),
    .X(_1417_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5314_ (.A0(rf_reg[413]),
    .A1(rf_reg[445]),
    .S(raddr_a_i[0]),
    .X(_1418_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5315_ (.Y(_1419_),
    .B1(_1418_),
    .B2(net259),
    .A2(_1417_),
    .A1(net275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5316_ (.A0(rf_reg[349]),
    .A1(rf_reg[381]),
    .S(raddr_a_i[0]),
    .X(_1420_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5317_ (.A0(rf_reg[285]),
    .A1(rf_reg[317]),
    .S(raddr_a_i[0]),
    .X(_1421_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5318_ (.Y(_1422_),
    .B1(_1421_),
    .B2(net248),
    .A2(_1420_),
    .A1(net237),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5319_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net232),
    .Y(_1423_),
    .A2(_1422_),
    .A1(_1419_));
 sg13g2_a221oi_1 _5320_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1423_),
    .B1(_1416_),
    .A1(net66),
    .Y(_1424_),
    .A2(_1415_));
 sg13g2_nand3_1 _5321_ (.B(_1414_),
    .C(_1424_),
    .A(_1405_),
    .Y(rdata_a_o[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5322_ (.A0(rf_reg[907]),
    .A1(rf_reg[939]),
    .S(raddr_a_i[0]),
    .X(_1425_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5323_ (.A0(rf_reg[971]),
    .A1(rf_reg[1003]),
    .S(raddr_a_i[0]),
    .X(_1426_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5324_ (.Y(_1427_),
    .B1(_1426_),
    .B2(net283),
    .A2(_1425_),
    .A1(net267),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(net266),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5326_ (.A0(rf_reg[779]),
    .A1(rf_reg[811]),
    .S(raddr_a_i[0]),
    .X(_1429_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5327_ (.A0(rf_reg[843]),
    .A1(rf_reg[875]),
    .S(raddr_a_i[0]),
    .X(_1430_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5328_ (.Y(_1431_),
    .B1(_1430_),
    .B2(net242),
    .A2(_1429_),
    .A1(net253),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 _5329_ (.A2(_1431_),
    .A1(_1427_),
    .B1(net309),
    .X(_1432_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5330_ (.A0(rf_reg[43]),
    .A1(rf_reg[107]),
    .S(raddr_a_i[1]),
    .X(_1433_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5331_ (.Y(_1434_),
    .A(raddr_a_i[0]),
    .B(_1433_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5332_ (.B(rf_reg[75]),
    .C(raddr_a_i[1]),
    .Y(_1435_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5333_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1434_),
    .A2(_1435_),
    .Y(_1436_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5334_ (.A0(rf_reg[139]),
    .A1(rf_reg[171]),
    .S(raddr_a_i[0]),
    .X(_1437_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5335_ (.A0(rf_reg[203]),
    .A1(rf_reg[235]),
    .S(raddr_a_i[0]),
    .X(_1438_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5336_ (.Y(_1439_),
    .B1(_1438_),
    .B2(net289),
    .A2(_1437_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5337_ (.VDD(VDD),
    .Y(_1440_),
    .A(_1439_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5338_ (.B1(net314),
    .VDD(VDD),
    .Y(_1441_),
    .VSS(VSS),
    .A1(_1436_),
    .A2(_1440_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5340_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[651]),
    .A1(rf_reg[683]),
    .A2(rf_reg[715]),
    .A3(rf_reg[747]),
    .S1(raddr_a_i[1]),
    .X(_1443_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5341_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[523]),
    .A1(rf_reg[555]),
    .A2(rf_reg[587]),
    .A3(rf_reg[619]),
    .S1(raddr_a_i[1]),
    .X(_1444_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5342_ (.A0(rf_reg[459]),
    .A1(rf_reg[491]),
    .S(raddr_a_i[0]),
    .X(_1445_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5343_ (.A0(rf_reg[395]),
    .A1(rf_reg[427]),
    .S(raddr_a_i[0]),
    .X(_1446_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5344_ (.Y(_1447_),
    .B1(_1446_),
    .B2(net267),
    .A2(_1445_),
    .A1(net283),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5345_ (.A0(rf_reg[331]),
    .A1(rf_reg[363]),
    .S(raddr_a_i[0]),
    .X(_1448_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5346_ (.A0(rf_reg[267]),
    .A1(rf_reg[299]),
    .S(raddr_a_i[0]),
    .X(_1449_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5347_ (.Y(_1450_),
    .B1(_1449_),
    .B2(net253),
    .A2(_1448_),
    .A1(net242),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5348_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net235),
    .Y(_1451_),
    .A2(_1450_),
    .A1(_1447_));
 sg13g2_a221oi_1 _5349_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1451_),
    .B1(_1444_),
    .A1(net69),
    .Y(_1452_),
    .A2(_1443_));
 sg13g2_nand3_1 _5350_ (.B(_1441_),
    .C(_1452_),
    .A(_1432_),
    .Y(rdata_a_o[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5351_ (.A0(rf_reg[906]),
    .A1(rf_reg[938]),
    .S(raddr_a_i[0]),
    .X(_1453_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5352_ (.A0(rf_reg[970]),
    .A1(rf_reg[1002]),
    .S(raddr_a_i[0]),
    .X(_1454_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5353_ (.Y(_1455_),
    .B1(_1454_),
    .B2(net278),
    .A2(_1453_),
    .A1(net262),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5354_ (.A0(rf_reg[778]),
    .A1(rf_reg[810]),
    .S(raddr_a_i[0]),
    .X(_1456_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5355_ (.A0(rf_reg[842]),
    .A1(rf_reg[874]),
    .S(raddr_a_i[0]),
    .X(_1457_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5356_ (.Y(_1458_),
    .B1(_1457_),
    .B2(net240),
    .A2(_1456_),
    .A1(net251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5357_ (.A2(_1458_),
    .A1(_1455_),
    .B1(net307),
    .X(_1459_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5358_ (.A0(rf_reg[42]),
    .A1(rf_reg[106]),
    .S(raddr_a_i[1]),
    .X(_1460_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5359_ (.Y(_1461_),
    .A(raddr_a_i[0]),
    .B(_1460_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5360_ (.B(rf_reg[74]),
    .C(raddr_a_i[1]),
    .Y(_1462_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5361_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1461_),
    .A2(_1462_),
    .Y(_1463_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5362_ (.A0(rf_reg[138]),
    .A1(rf_reg[170]),
    .S(raddr_a_i[0]),
    .X(_1464_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5363_ (.A0(rf_reg[202]),
    .A1(rf_reg[234]),
    .S(raddr_a_i[0]),
    .X(_1465_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5364_ (.Y(_1466_),
    .B1(_1465_),
    .B2(net281),
    .A2(_1464_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5365_ (.VDD(VDD),
    .Y(_1467_),
    .A(_1466_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5366_ (.B1(net312),
    .VDD(VDD),
    .Y(_1468_),
    .VSS(VSS),
    .A1(_1463_),
    .A2(_1467_));
 sg13g2_mux4_1 _5367_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[650]),
    .A1(rf_reg[682]),
    .A2(rf_reg[714]),
    .A3(rf_reg[746]),
    .S1(raddr_a_i[1]),
    .X(_1469_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5368_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[522]),
    .A1(rf_reg[554]),
    .A2(rf_reg[586]),
    .A3(rf_reg[618]),
    .S1(raddr_a_i[1]),
    .X(_1470_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5369_ (.A0(rf_reg[458]),
    .A1(rf_reg[490]),
    .S(raddr_a_i[0]),
    .X(_1471_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5370_ (.A0(rf_reg[394]),
    .A1(rf_reg[426]),
    .S(raddr_a_i[0]),
    .X(_1472_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5371_ (.Y(_1473_),
    .B1(_1472_),
    .B2(net261),
    .A2(_1471_),
    .A1(net277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5372_ (.A0(rf_reg[330]),
    .A1(rf_reg[362]),
    .S(raddr_a_i[0]),
    .X(_1474_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5373_ (.A0(rf_reg[266]),
    .A1(rf_reg[298]),
    .S(raddr_a_i[0]),
    .X(_1475_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5374_ (.Y(_1476_),
    .B1(_1475_),
    .B2(net250),
    .A2(_1474_),
    .A1(net239),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5375_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net233),
    .Y(_1477_),
    .A2(_1476_),
    .A1(_1473_));
 sg13g2_a221oi_1 _5376_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net228),
    .C1(_1477_),
    .B1(_1470_),
    .A1(net67),
    .Y(_1478_),
    .A2(_1469_));
 sg13g2_nand3_1 _5377_ (.B(_1468_),
    .C(_1478_),
    .A(_1459_),
    .Y(rdata_a_o[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5378_ (.A0(rf_reg[905]),
    .A1(rf_reg[937]),
    .S(raddr_a_i[0]),
    .X(_1479_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5379_ (.A0(rf_reg[969]),
    .A1(rf_reg[1001]),
    .S(raddr_a_i[0]),
    .X(_1480_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5380_ (.Y(_1481_),
    .B1(_1480_),
    .B2(net275),
    .A2(_1479_),
    .A1(net259),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5381_ (.A0(rf_reg[777]),
    .A1(rf_reg[809]),
    .S(raddr_a_i[0]),
    .X(_1482_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5382_ (.A0(rf_reg[841]),
    .A1(rf_reg[873]),
    .S(raddr_a_i[0]),
    .X(_1483_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5383_ (.Y(_1484_),
    .B1(_1483_),
    .B2(net238),
    .A2(_1482_),
    .A1(net249),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5384_ (.A2(_1484_),
    .A1(_1481_),
    .B1(net306),
    .X(_1485_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net266),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5386_ (.A0(rf_reg[41]),
    .A1(rf_reg[105]),
    .S(raddr_a_i[1]),
    .X(_1487_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5387_ (.Y(_1488_),
    .A(raddr_a_i[0]),
    .B(_1487_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5388_ (.B(rf_reg[73]),
    .C(raddr_a_i[1]),
    .Y(_1489_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5389_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1488_),
    .A2(_1489_),
    .Y(_1490_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5390_ (.A0(rf_reg[137]),
    .A1(rf_reg[169]),
    .S(raddr_a_i[0]),
    .X(_1491_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5391_ (.A0(rf_reg[201]),
    .A1(rf_reg[233]),
    .S(raddr_a_i[0]),
    .X(_1492_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5392_ (.Y(_1493_),
    .B1(_1492_),
    .B2(net280),
    .A2(_1491_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5393_ (.VDD(VDD),
    .Y(_1494_),
    .A(_1493_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5394_ (.B1(net311),
    .VDD(VDD),
    .Y(_1495_),
    .VSS(VSS),
    .A1(_1490_),
    .A2(_1494_));
 sg13g2_mux4_1 _5395_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[649]),
    .A1(rf_reg[681]),
    .A2(rf_reg[713]),
    .A3(rf_reg[745]),
    .S1(raddr_a_i[1]),
    .X(_1496_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5396_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[521]),
    .A1(rf_reg[553]),
    .A2(rf_reg[585]),
    .A3(rf_reg[617]),
    .S1(raddr_a_i[1]),
    .X(_1497_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5397_ (.A0(rf_reg[457]),
    .A1(rf_reg[489]),
    .S(raddr_a_i[0]),
    .X(_1498_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5398_ (.A0(rf_reg[393]),
    .A1(rf_reg[425]),
    .S(raddr_a_i[0]),
    .X(_1499_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5399_ (.Y(_1500_),
    .B1(_1499_),
    .B2(net259),
    .A2(_1498_),
    .A1(net275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5400_ (.A0(rf_reg[329]),
    .A1(rf_reg[361]),
    .S(raddr_a_i[0]),
    .X(_1501_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(net263),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5402_ (.A0(rf_reg[265]),
    .A1(rf_reg[297]),
    .S(raddr_a_i[0]),
    .X(_1503_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5403_ (.Y(_1504_),
    .B1(_1503_),
    .B2(net249),
    .A2(_1501_),
    .A1(net238),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5404_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net232),
    .Y(_1505_),
    .A2(_1504_),
    .A1(_1500_));
 sg13g2_a221oi_1 _5405_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1505_),
    .B1(_1497_),
    .A1(net66),
    .Y(_1506_),
    .A2(_1496_));
 sg13g2_nand3_1 _5406_ (.B(_1495_),
    .C(_1506_),
    .A(_1485_),
    .Y(rdata_a_o[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5407_ (.A0(rf_reg[904]),
    .A1(rf_reg[936]),
    .S(raddr_a_i[0]),
    .X(_1507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5408_ (.A0(rf_reg[968]),
    .A1(rf_reg[1000]),
    .S(raddr_a_i[0]),
    .X(_1508_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5409_ (.Y(_1509_),
    .B1(_1508_),
    .B2(net277),
    .A2(_1507_),
    .A1(net261),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5410_ (.A0(rf_reg[776]),
    .A1(rf_reg[808]),
    .S(raddr_a_i[0]),
    .X(_1510_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5411_ (.A0(rf_reg[840]),
    .A1(rf_reg[872]),
    .S(raddr_a_i[0]),
    .X(_1511_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5412_ (.Y(_1512_),
    .B1(_1511_),
    .B2(net239),
    .A2(_1510_),
    .A1(net250),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5413_ (.A2(_1512_),
    .A1(_1509_),
    .B1(net306),
    .X(_1513_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5414_ (.A0(rf_reg[40]),
    .A1(rf_reg[104]),
    .S(raddr_a_i[1]),
    .X(_1514_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5415_ (.Y(_1515_),
    .A(raddr_a_i[0]),
    .B(_1514_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net262),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5417_ (.B(rf_reg[72]),
    .C(raddr_a_i[1]),
    .Y(_1517_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5418_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1515_),
    .A2(_1517_),
    .Y(_1518_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5419_ (.A0(rf_reg[136]),
    .A1(rf_reg[168]),
    .S(raddr_a_i[0]),
    .X(_1519_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5420_ (.A0(rf_reg[200]),
    .A1(rf_reg[232]),
    .S(raddr_a_i[0]),
    .X(_1520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5421_ (.Y(_1521_),
    .B1(_1520_),
    .B2(net280),
    .A2(_1519_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5422_ (.VDD(VDD),
    .Y(_1522_),
    .A(_1521_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5423_ (.B1(net312),
    .VDD(VDD),
    .Y(_1523_),
    .VSS(VSS),
    .A1(_1518_),
    .A2(_1522_));
 sg13g2_mux4_1 _5424_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[648]),
    .A1(rf_reg[680]),
    .A2(rf_reg[712]),
    .A3(rf_reg[744]),
    .S1(raddr_a_i[1]),
    .X(_1524_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5425_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[520]),
    .A1(rf_reg[552]),
    .A2(rf_reg[584]),
    .A3(rf_reg[616]),
    .S1(raddr_a_i[1]),
    .X(_1525_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(net263),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5427_ (.A0(rf_reg[456]),
    .A1(rf_reg[488]),
    .S(raddr_a_i[0]),
    .X(_1527_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5428_ (.A0(rf_reg[392]),
    .A1(rf_reg[424]),
    .S(raddr_a_i[0]),
    .X(_1528_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(net263),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5430_ (.Y(_1530_),
    .B1(_1528_),
    .B2(net261),
    .A2(_1527_),
    .A1(net277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5431_ (.A0(rf_reg[328]),
    .A1(rf_reg[360]),
    .S(raddr_a_i[0]),
    .X(_1531_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5432_ (.A0(rf_reg[264]),
    .A1(rf_reg[296]),
    .S(raddr_a_i[0]),
    .X(_1532_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5433_ (.Y(_1533_),
    .B1(_1532_),
    .B2(net250),
    .A2(_1531_),
    .A1(net239),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5434_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net233),
    .Y(_1534_),
    .A2(_1533_),
    .A1(_1530_));
 sg13g2_a221oi_1 _5435_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1534_),
    .B1(_1525_),
    .A1(net66),
    .Y(_1535_),
    .A2(_1524_));
 sg13g2_nand3_1 _5436_ (.B(_1523_),
    .C(_1535_),
    .A(_1513_),
    .Y(rdata_a_o[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout258 (.A(_1010_),
    .X(net258),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5438_ (.A0(rf_reg[903]),
    .A1(rf_reg[935]),
    .S(raddr_a_i[0]),
    .X(_1537_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5439_ (.A0(rf_reg[967]),
    .A1(rf_reg[999]),
    .S(raddr_a_i[0]),
    .X(_1538_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5440_ (.Y(_1539_),
    .B1(_1538_),
    .B2(net288),
    .A2(_1537_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5441_ (.A0(rf_reg[775]),
    .A1(rf_reg[807]),
    .S(raddr_a_i[0]),
    .X(_1540_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5442_ (.A0(rf_reg[839]),
    .A1(rf_reg[871]),
    .S(raddr_a_i[0]),
    .X(_1541_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5443_ (.Y(_1542_),
    .B1(_1541_),
    .B2(net245),
    .A2(_1540_),
    .A1(net256),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5444_ (.A2(_1542_),
    .A1(_1539_),
    .B1(net308),
    .X(_1543_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5445_ (.A0(rf_reg[39]),
    .A1(rf_reg[103]),
    .S(raddr_a_i[1]),
    .X(_1544_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5446_ (.Y(_1545_),
    .A(raddr_a_i[0]),
    .B(_1544_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5447_ (.B(rf_reg[71]),
    .C(raddr_a_i[1]),
    .Y(_1546_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5448_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1545_),
    .A2(_1546_),
    .Y(_1547_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5449_ (.A0(rf_reg[135]),
    .A1(rf_reg[167]),
    .S(raddr_a_i[0]),
    .X(_1548_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5450_ (.A0(rf_reg[199]),
    .A1(rf_reg[231]),
    .S(raddr_a_i[0]),
    .X(_1549_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5451_ (.Y(_1550_),
    .B1(_1549_),
    .B2(net288),
    .A2(_1548_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5452_ (.VDD(VDD),
    .Y(_1551_),
    .A(_1550_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5453_ (.B1(net313),
    .VDD(VDD),
    .Y(_1552_),
    .VSS(VSS),
    .A1(_1547_),
    .A2(_1551_));
 sg13g2_mux4_1 _5454_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[647]),
    .A1(rf_reg[679]),
    .A2(rf_reg[711]),
    .A3(rf_reg[743]),
    .S1(raddr_a_i[1]),
    .X(_1553_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5456_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[519]),
    .A1(rf_reg[551]),
    .A2(rf_reg[583]),
    .A3(rf_reg[615]),
    .S1(raddr_a_i[1]),
    .X(_1555_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5457_ (.A0(rf_reg[455]),
    .A1(rf_reg[487]),
    .S(raddr_a_i[0]),
    .X(_1556_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(net257),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5459_ (.A0(rf_reg[391]),
    .A1(rf_reg[423]),
    .S(raddr_a_i[0]),
    .X(_1558_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5460_ (.Y(_1559_),
    .B1(_1558_),
    .B2(net270),
    .A2(_1556_),
    .A1(net286),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5461_ (.A0(rf_reg[327]),
    .A1(rf_reg[359]),
    .S(raddr_a_i[0]),
    .X(_1560_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5462_ (.A0(rf_reg[263]),
    .A1(rf_reg[295]),
    .S(raddr_a_i[0]),
    .X(_1561_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5463_ (.Y(_1562_),
    .B1(_1561_),
    .B2(net256),
    .A2(_1560_),
    .A1(net245),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5464_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1559_),
    .A2(_1562_),
    .Y(_1563_),
    .B1(net234));
 sg13g2_a221oi_1 _5465_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1563_),
    .B1(_1555_),
    .A1(net68),
    .Y(_1564_),
    .A2(_1553_));
 sg13g2_nand3_1 _5466_ (.B(_1552_),
    .C(_1564_),
    .A(_1543_),
    .Y(rdata_a_o[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5467_ (.A0(rf_reg[902]),
    .A1(rf_reg[934]),
    .S(raddr_a_i[0]),
    .X(_1565_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5468_ (.A0(rf_reg[966]),
    .A1(rf_reg[998]),
    .S(raddr_a_i[0]),
    .X(_1566_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5469_ (.Y(_1567_),
    .B1(_1566_),
    .B2(net278),
    .A2(_1565_),
    .A1(net262),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5470_ (.A0(rf_reg[774]),
    .A1(rf_reg[806]),
    .S(raddr_a_i[0]),
    .X(_1568_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5471_ (.A0(rf_reg[838]),
    .A1(rf_reg[870]),
    .S(raddr_a_i[0]),
    .X(_1569_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5472_ (.Y(_1570_),
    .B1(_1569_),
    .B2(net240),
    .A2(_1568_),
    .A1(net251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5473_ (.A2(_1570_),
    .A1(_1567_),
    .B1(net307),
    .X(_1571_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5474_ (.A0(rf_reg[38]),
    .A1(rf_reg[102]),
    .S(raddr_a_i[1]),
    .X(_1572_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5475_ (.Y(_1573_),
    .A(raddr_a_i[0]),
    .B(_1572_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(net257),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5477_ (.B(rf_reg[70]),
    .C(raddr_a_i[1]),
    .Y(_1575_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5478_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1573_),
    .A2(_1575_),
    .Y(_1576_),
    .B1(raddr_a_i[2]));
 sg13g2_buf_2 fanout254 (.A(net258),
    .X(net254),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5480_ (.A0(rf_reg[134]),
    .A1(rf_reg[166]),
    .S(raddr_a_i[0]),
    .X(_1578_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5481_ (.A0(rf_reg[198]),
    .A1(rf_reg[230]),
    .S(raddr_a_i[0]),
    .X(_1579_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(net258),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5483_ (.Y(_1581_),
    .B1(_1579_),
    .B2(net282),
    .A2(_1578_),
    .A1(net266),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5484_ (.VDD(VDD),
    .Y(_1582_),
    .A(_1581_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5485_ (.B1(net311),
    .VDD(VDD),
    .Y(_1583_),
    .VSS(VSS),
    .A1(_1576_),
    .A2(_1582_));
 sg13g2_buf_2 fanout252 (.A(net258),
    .X(net252),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5487_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[646]),
    .A1(rf_reg[678]),
    .A2(rf_reg[710]),
    .A3(rf_reg[742]),
    .S1(raddr_a_i[1]),
    .X(_1585_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5488_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[518]),
    .A1(rf_reg[550]),
    .A2(rf_reg[582]),
    .A3(rf_reg[614]),
    .S1(raddr_a_i[1]),
    .X(_1586_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5489_ (.A0(rf_reg[454]),
    .A1(rf_reg[486]),
    .S(raddr_a_i[0]),
    .X(_1587_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5490_ (.A0(rf_reg[390]),
    .A1(rf_reg[422]),
    .S(raddr_a_i[0]),
    .X(_1588_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5491_ (.Y(_1589_),
    .B1(_1588_),
    .B2(net263),
    .A2(_1587_),
    .A1(net278),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(net252),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(net251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5494_ (.A0(rf_reg[326]),
    .A1(rf_reg[358]),
    .S(raddr_a_i[0]),
    .X(_1592_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5495_ (.A0(rf_reg[262]),
    .A1(rf_reg[294]),
    .S(raddr_a_i[0]),
    .X(_1593_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(net252),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5497_ (.Y(_1595_),
    .B1(_1593_),
    .B2(net252),
    .A2(_1592_),
    .A1(net241),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5498_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net233),
    .Y(_1596_),
    .A2(_1595_),
    .A1(_1589_));
 sg13g2_a221oi_1 _5499_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net228),
    .C1(_1596_),
    .B1(_1586_),
    .A1(net67),
    .Y(_1597_),
    .A2(_1585_));
 sg13g2_nand3_1 _5500_ (.B(_1583_),
    .C(_1597_),
    .A(_1571_),
    .Y(rdata_a_o[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5501_ (.A0(rf_reg[901]),
    .A1(rf_reg[933]),
    .S(raddr_a_i[0]),
    .X(_1598_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5502_ (.A0(rf_reg[965]),
    .A1(rf_reg[997]),
    .S(raddr_a_i[0]),
    .X(_1599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5503_ (.Y(_1600_),
    .B1(_1599_),
    .B2(net285),
    .A2(_1598_),
    .A1(net269),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5504_ (.A0(rf_reg[773]),
    .A1(rf_reg[805]),
    .S(raddr_a_i[0]),
    .X(_1601_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5505_ (.A0(rf_reg[837]),
    .A1(rf_reg[869]),
    .S(raddr_a_i[0]),
    .X(_1602_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5506_ (.Y(_1603_),
    .B1(_1602_),
    .B2(net245),
    .A2(_1601_),
    .A1(net256),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5507_ (.A2(_1603_),
    .A1(_1600_),
    .B1(net308),
    .X(_1604_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5508_ (.A0(rf_reg[37]),
    .A1(rf_reg[101]),
    .S(raddr_a_i[1]),
    .X(_1605_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5509_ (.Y(_1606_),
    .A(raddr_a_i[0]),
    .B(_1605_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5510_ (.B(rf_reg[69]),
    .C(raddr_a_i[1]),
    .Y(_1607_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5511_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1606_),
    .A2(_1607_),
    .Y(_1608_),
    .B1(raddr_a_i[2]));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net249),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5513_ (.A0(rf_reg[133]),
    .A1(rf_reg[165]),
    .S(raddr_a_i[0]),
    .X(_1610_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5514_ (.A0(rf_reg[197]),
    .A1(rf_reg[229]),
    .S(raddr_a_i[0]),
    .X(_1611_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5515_ (.Y(_1612_),
    .B1(_1611_),
    .B2(net290),
    .A2(_1610_),
    .A1(net274),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5516_ (.VDD(VDD),
    .Y(_1613_),
    .A(_1612_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5517_ (.B1(net313),
    .VDD(VDD),
    .Y(_1614_),
    .VSS(VSS),
    .A1(_1608_),
    .A2(_1613_));
 sg13g2_mux4_1 _5518_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[645]),
    .A1(rf_reg[677]),
    .A2(rf_reg[709]),
    .A3(rf_reg[741]),
    .S1(raddr_a_i[1]),
    .X(_1615_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5519_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[517]),
    .A1(rf_reg[549]),
    .A2(rf_reg[581]),
    .A3(rf_reg[613]),
    .S1(raddr_a_i[1]),
    .X(_1616_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5520_ (.A0(rf_reg[453]),
    .A1(rf_reg[485]),
    .S(raddr_a_i[0]),
    .X(_1617_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5521_ (.A0(rf_reg[389]),
    .A1(rf_reg[421]),
    .S(raddr_a_i[0]),
    .X(_1618_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5522_ (.Y(_1619_),
    .B1(_1618_),
    .B2(net270),
    .A2(_1617_),
    .A1(net286),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5523_ (.A0(rf_reg[325]),
    .A1(rf_reg[357]),
    .S(raddr_a_i[0]),
    .X(_1620_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5524_ (.A0(rf_reg[261]),
    .A1(rf_reg[293]),
    .S(raddr_a_i[0]),
    .X(_1621_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5525_ (.Y(_1622_),
    .B1(_1621_),
    .B2(net256),
    .A2(_1620_),
    .A1(net246),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5526_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1619_),
    .A2(_1622_),
    .Y(_1623_),
    .B1(net234));
 sg13g2_a221oi_1 _5527_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1623_),
    .B1(_1616_),
    .A1(net68),
    .Y(_1624_),
    .A2(_1615_));
 sg13g2_nand3_1 _5528_ (.B(_1614_),
    .C(_1624_),
    .A(_1604_),
    .Y(rdata_a_o[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout247 (.A(_1014_),
    .X(net247),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5530_ (.A0(rf_reg[900]),
    .A1(rf_reg[932]),
    .S(raddr_a_i[0]),
    .X(_1626_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5531_ (.A0(rf_reg[964]),
    .A1(rf_reg[996]),
    .S(raddr_a_i[0]),
    .X(_1627_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5532_ (.Y(_1628_),
    .B1(_1627_),
    .B2(net276),
    .A2(_1626_),
    .A1(net260),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5533_ (.A0(rf_reg[772]),
    .A1(rf_reg[804]),
    .S(raddr_a_i[0]),
    .X(_1629_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(net247),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5535_ (.A0(rf_reg[836]),
    .A1(rf_reg[868]),
    .S(raddr_a_i[0]),
    .X(_1631_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(net246),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5537_ (.Y(_1633_),
    .B1(_1631_),
    .B2(net241),
    .A2(_1629_),
    .A1(net252),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5538_ (.A2(_1633_),
    .A1(_1628_),
    .B1(net306),
    .X(_1634_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(net246),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5540_ (.A0(rf_reg[36]),
    .A1(rf_reg[100]),
    .S(raddr_a_i[1]),
    .X(_1636_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5541_ (.Y(_1637_),
    .A(raddr_a_i[0]),
    .B(_1636_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5542_ (.B(rf_reg[68]),
    .C(raddr_a_i[1]),
    .Y(_1638_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_buf_2 fanout243 (.A(net247),
    .X(net243),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5544_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1637_),
    .A2(_1638_),
    .Y(_1640_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5545_ (.A0(rf_reg[132]),
    .A1(rf_reg[164]),
    .S(raddr_a_i[0]),
    .X(_1641_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5546_ (.A0(rf_reg[196]),
    .A1(rf_reg[228]),
    .S(raddr_a_i[0]),
    .X(_1642_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5547_ (.Y(_1643_),
    .B1(_1642_),
    .B2(net280),
    .A2(_1641_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5548_ (.VDD(VDD),
    .Y(_1644_),
    .A(_1643_),
    .VSS(VSS));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(net247),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _5550_ (.B1(net311),
    .VDD(VDD),
    .Y(_1646_),
    .VSS(VSS),
    .A1(_1640_),
    .A2(_1644_));
 sg13g2_buf_2 fanout241 (.A(net247),
    .X(net241),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5552_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[644]),
    .A1(rf_reg[676]),
    .A2(rf_reg[708]),
    .A3(rf_reg[740]),
    .S1(raddr_a_i[1]),
    .X(_1648_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5553_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[516]),
    .A1(rf_reg[548]),
    .A2(rf_reg[580]),
    .A3(rf_reg[612]),
    .S1(raddr_a_i[1]),
    .X(_1649_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(net241),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(net240),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5556_ (.A0(rf_reg[452]),
    .A1(rf_reg[484]),
    .S(raddr_a_i[0]),
    .X(_1652_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5557_ (.A0(rf_reg[388]),
    .A1(rf_reg[420]),
    .S(raddr_a_i[0]),
    .X(_1653_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5558_ (.Y(_1654_),
    .B1(_1653_),
    .B2(net259),
    .A2(_1652_),
    .A1(net275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5559_ (.A0(rf_reg[324]),
    .A1(rf_reg[356]),
    .S(raddr_a_i[0]),
    .X(_1655_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5560_ (.A0(rf_reg[260]),
    .A1(rf_reg[292]),
    .S(raddr_a_i[0]),
    .X(_1656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5561_ (.Y(_1657_),
    .B1(_1656_),
    .B2(net249),
    .A2(_1655_),
    .A1(net238),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(net241),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5563_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net232),
    .Y(_1659_),
    .A2(_1657_),
    .A1(_1654_));
 sg13g2_a221oi_1 _5564_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net228),
    .C1(_1659_),
    .B1(_1649_),
    .A1(net67),
    .Y(_1660_),
    .A2(_1648_));
 sg13g2_nand3_1 _5565_ (.B(_1646_),
    .C(_1660_),
    .A(_1634_),
    .Y(rdata_a_o[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5566_ (.A0(rf_reg[899]),
    .A1(rf_reg[931]),
    .S(raddr_a_i[0]),
    .X(_1661_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5567_ (.A0(rf_reg[963]),
    .A1(rf_reg[995]),
    .S(raddr_a_i[0]),
    .X(_1662_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(net238),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5569_ (.Y(_1664_),
    .B1(_1662_),
    .B2(net287),
    .A2(_1661_),
    .A1(net271),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(_1019_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5571_ (.A0(rf_reg[771]),
    .A1(rf_reg[803]),
    .S(raddr_a_i[0]),
    .X(_1666_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5572_ (.A0(rf_reg[835]),
    .A1(rf_reg[867]),
    .S(raddr_a_i[0]),
    .X(_1667_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5573_ (.Y(_1668_),
    .B1(_1667_),
    .B2(net246),
    .A2(_1666_),
    .A1(net257),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(net236),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5575_ (.A2(_1668_),
    .A1(_1664_),
    .B1(net309),
    .X(_1670_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5576_ (.A0(rf_reg[35]),
    .A1(rf_reg[99]),
    .S(raddr_a_i[1]),
    .X(_1671_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5577_ (.Y(_1672_),
    .A(raddr_a_i[0]),
    .B(_1671_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5578_ (.B(rf_reg[67]),
    .C(raddr_a_i[1]),
    .Y(_1673_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5579_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1672_),
    .A2(_1673_),
    .Y(_1674_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5580_ (.A0(rf_reg[131]),
    .A1(rf_reg[163]),
    .S(raddr_a_i[0]),
    .X(_1675_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(net235),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5582_ (.A0(rf_reg[195]),
    .A1(rf_reg[227]),
    .S(raddr_a_i[0]),
    .X(_1677_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5583_ (.Y(_1678_),
    .B1(_1677_),
    .B2(net288),
    .A2(_1675_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5584_ (.VDD(VDD),
    .Y(_1679_),
    .A(_1678_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5585_ (.B1(net314),
    .VDD(VDD),
    .Y(_1680_),
    .VSS(VSS),
    .A1(_1674_),
    .A2(_1679_));
 sg13g2_mux4_1 _5586_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[643]),
    .A1(rf_reg[675]),
    .A2(rf_reg[707]),
    .A3(rf_reg[739]),
    .S1(raddr_a_i[1]),
    .X(_1681_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(net236),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5588_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[515]),
    .A1(rf_reg[547]),
    .A2(rf_reg[579]),
    .A3(rf_reg[611]),
    .S1(raddr_a_i[1]),
    .X(_1683_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5589_ (.A0(rf_reg[451]),
    .A1(rf_reg[483]),
    .S(raddr_a_i[0]),
    .X(_1684_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5590_ (.A0(rf_reg[387]),
    .A1(rf_reg[419]),
    .S(raddr_a_i[0]),
    .X(_1685_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5591_ (.Y(_1686_),
    .B1(_1685_),
    .B2(net270),
    .A2(_1684_),
    .A1(net286),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5592_ (.A0(rf_reg[323]),
    .A1(rf_reg[355]),
    .S(raddr_a_i[0]),
    .X(_1687_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5593_ (.A0(rf_reg[259]),
    .A1(rf_reg[291]),
    .S(raddr_a_i[0]),
    .X(_1688_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5594_ (.Y(_1689_),
    .B1(_1688_),
    .B2(net256),
    .A2(_1687_),
    .A1(net245),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5595_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1686_),
    .A2(_1689_),
    .Y(_1690_),
    .B1(net235));
 sg13g2_a221oi_1 _5596_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1690_),
    .B1(_1683_),
    .A1(net69),
    .Y(_1691_),
    .A2(_1681_));
 sg13g2_nand3_1 _5597_ (.B(_1680_),
    .C(_1691_),
    .A(_1670_),
    .Y(rdata_a_o[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5598_ (.A0(rf_reg[898]),
    .A1(rf_reg[930]),
    .S(raddr_a_i[0]),
    .X(_1692_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(net236),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5600_ (.A0(rf_reg[962]),
    .A1(rf_reg[994]),
    .S(raddr_a_i[0]),
    .X(_1694_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5601_ (.Y(_1695_),
    .B1(_1694_),
    .B2(net275),
    .A2(_1692_),
    .A1(net259),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5602_ (.A0(rf_reg[770]),
    .A1(rf_reg[802]),
    .S(raddr_a_i[0]),
    .X(_1696_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5603_ (.A0(rf_reg[834]),
    .A1(rf_reg[866]),
    .S(raddr_a_i[0]),
    .X(_1697_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5604_ (.Y(_1698_),
    .B1(_1697_),
    .B2(net238),
    .A2(_1696_),
    .A1(net249),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5605_ (.A2(_1698_),
    .A1(_1695_),
    .B1(net306),
    .X(_1699_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5606_ (.A0(rf_reg[34]),
    .A1(rf_reg[98]),
    .S(raddr_a_i[1]),
    .X(_1700_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5607_ (.Y(_1701_),
    .A(raddr_a_i[0]),
    .B(_1700_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5608_ (.B(rf_reg[66]),
    .C(raddr_a_i[1]),
    .Y(_1702_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5609_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1701_),
    .A2(_1702_),
    .Y(_1703_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5610_ (.A0(rf_reg[130]),
    .A1(rf_reg[162]),
    .S(raddr_a_i[0]),
    .X(_1704_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5611_ (.A0(rf_reg[194]),
    .A1(rf_reg[226]),
    .S(raddr_a_i[0]),
    .X(_1705_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5612_ (.Y(_1706_),
    .B1(_1705_),
    .B2(net281),
    .A2(_1704_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5613_ (.VDD(VDD),
    .Y(_1707_),
    .A(_1706_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5614_ (.B1(net311),
    .VDD(VDD),
    .Y(_1708_),
    .VSS(VSS),
    .A1(_1703_),
    .A2(_1707_));
 sg13g2_mux4_1 _5615_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[642]),
    .A1(rf_reg[674]),
    .A2(rf_reg[706]),
    .A3(rf_reg[738]),
    .S1(raddr_a_i[1]),
    .X(_1709_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5616_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[514]),
    .A1(rf_reg[546]),
    .A2(rf_reg[578]),
    .A3(rf_reg[610]),
    .S1(raddr_a_i[1]),
    .X(_1710_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5617_ (.A0(rf_reg[450]),
    .A1(rf_reg[482]),
    .S(raddr_a_i[0]),
    .X(_1711_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5618_ (.A0(rf_reg[386]),
    .A1(rf_reg[418]),
    .S(raddr_a_i[0]),
    .X(_1712_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5619_ (.Y(_1713_),
    .B1(_1712_),
    .B2(net259),
    .A2(_1711_),
    .A1(net275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5620_ (.A0(rf_reg[322]),
    .A1(rf_reg[354]),
    .S(raddr_a_i[0]),
    .X(_1714_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5621_ (.A0(rf_reg[258]),
    .A1(rf_reg[290]),
    .S(raddr_a_i[0]),
    .X(_1715_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5622_ (.Y(_1716_),
    .B1(_1715_),
    .B2(net249),
    .A2(_1714_),
    .A1(net238),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5623_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net232),
    .Y(_1717_),
    .A2(_1716_),
    .A1(_1713_));
 sg13g2_a221oi_1 _5624_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1717_),
    .B1(_1710_),
    .A1(net66),
    .Y(_1718_),
    .A2(_1709_));
 sg13g2_nand3_1 _5625_ (.B(_1708_),
    .C(_1718_),
    .A(_1699_),
    .Y(rdata_a_o[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5626_ (.A0(rf_reg[924]),
    .A1(rf_reg[956]),
    .S(raddr_a_i[0]),
    .X(_1719_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5627_ (.A0(rf_reg[988]),
    .A1(rf_reg[1020]),
    .S(raddr_a_i[0]),
    .X(_1720_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5628_ (.Y(_1721_),
    .B1(_1720_),
    .B2(net286),
    .A2(_1719_),
    .A1(net270),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5629_ (.A0(rf_reg[796]),
    .A1(rf_reg[828]),
    .S(raddr_a_i[0]),
    .X(_1722_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5630_ (.A0(rf_reg[860]),
    .A1(rf_reg[892]),
    .S(raddr_a_i[0]),
    .X(_1723_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5631_ (.Y(_1724_),
    .B1(_1723_),
    .B2(net246),
    .A2(_1722_),
    .A1(net257),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5632_ (.A2(_1724_),
    .A1(_1721_),
    .B1(net308),
    .X(_1725_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5633_ (.A0(rf_reg[60]),
    .A1(rf_reg[124]),
    .S(raddr_a_i[1]),
    .X(_1726_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5634_ (.Y(_1727_),
    .A(raddr_a_i[0]),
    .B(_1726_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5635_ (.B(rf_reg[92]),
    .C(raddr_a_i[1]),
    .Y(_1728_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5636_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1727_),
    .A2(_1728_),
    .Y(_1729_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5637_ (.A0(rf_reg[156]),
    .A1(rf_reg[188]),
    .S(raddr_a_i[0]),
    .X(_1730_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5638_ (.A0(rf_reg[220]),
    .A1(rf_reg[252]),
    .S(raddr_a_i[0]),
    .X(_1731_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5639_ (.Y(_1732_),
    .B1(_1731_),
    .B2(net288),
    .A2(_1730_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5640_ (.VDD(VDD),
    .Y(_1733_),
    .A(_1732_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5641_ (.B1(net314),
    .VDD(VDD),
    .Y(_1734_),
    .VSS(VSS),
    .A1(_1729_),
    .A2(_1733_));
 sg13g2_mux4_1 _5642_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[668]),
    .A1(rf_reg[700]),
    .A2(rf_reg[732]),
    .A3(rf_reg[764]),
    .S1(raddr_a_i[1]),
    .X(_1735_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5643_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[540]),
    .A1(rf_reg[572]),
    .A2(rf_reg[604]),
    .A3(rf_reg[636]),
    .S1(raddr_a_i[1]),
    .X(_1736_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5644_ (.A0(rf_reg[476]),
    .A1(rf_reg[508]),
    .S(raddr_a_i[0]),
    .X(_1737_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5645_ (.A0(rf_reg[412]),
    .A1(rf_reg[444]),
    .S(raddr_a_i[0]),
    .X(_1738_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5646_ (.Y(_1739_),
    .B1(_1738_),
    .B2(net269),
    .A2(_1737_),
    .A1(net285),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5647_ (.A0(rf_reg[348]),
    .A1(rf_reg[380]),
    .S(raddr_a_i[0]),
    .X(_1740_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5648_ (.A0(rf_reg[284]),
    .A1(rf_reg[316]),
    .S(raddr_a_i[0]),
    .X(_1741_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5649_ (.Y(_1742_),
    .B1(_1741_),
    .B2(net255),
    .A2(_1740_),
    .A1(net246),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5650_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net234),
    .Y(_1743_),
    .A2(_1742_),
    .A1(_1739_));
 sg13g2_a221oi_1 _5651_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1743_),
    .B1(_1736_),
    .A1(net69),
    .Y(_1744_),
    .A2(_1735_));
 sg13g2_nand3_1 _5652_ (.B(_1734_),
    .C(_1744_),
    .A(_1725_),
    .Y(rdata_a_o[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5653_ (.A0(rf_reg[897]),
    .A1(rf_reg[929]),
    .S(raddr_a_i[0]),
    .X(_1745_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5654_ (.A0(rf_reg[961]),
    .A1(rf_reg[993]),
    .S(raddr_a_i[0]),
    .X(_1746_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5655_ (.Y(_1747_),
    .B1(_1746_),
    .B2(net283),
    .A2(_1745_),
    .A1(net267),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5656_ (.A0(rf_reg[769]),
    .A1(rf_reg[801]),
    .S(raddr_a_i[0]),
    .X(_1748_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5657_ (.A0(rf_reg[833]),
    .A1(rf_reg[865]),
    .S(raddr_a_i[0]),
    .X(_1749_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5658_ (.Y(_1750_),
    .B1(_1749_),
    .B2(net242),
    .A2(_1748_),
    .A1(net253),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5659_ (.A2(_1750_),
    .A1(_1747_),
    .B1(net309),
    .X(_1751_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5660_ (.A0(rf_reg[33]),
    .A1(rf_reg[97]),
    .S(raddr_a_i[1]),
    .X(_1752_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5661_ (.Y(_1753_),
    .A(raddr_a_i[0]),
    .B(_1752_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5662_ (.B(rf_reg[65]),
    .C(raddr_a_i[1]),
    .Y(_1754_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5663_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1753_),
    .A2(_1754_),
    .Y(_1755_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5664_ (.A0(rf_reg[129]),
    .A1(rf_reg[161]),
    .S(raddr_a_i[0]),
    .X(_1756_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5665_ (.A0(rf_reg[193]),
    .A1(rf_reg[225]),
    .S(raddr_a_i[0]),
    .X(_1757_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5666_ (.Y(_1758_),
    .B1(_1757_),
    .B2(net289),
    .A2(_1756_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5667_ (.VDD(VDD),
    .Y(_1759_),
    .A(_1758_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5668_ (.B1(net314),
    .VDD(VDD),
    .Y(_1760_),
    .VSS(VSS),
    .A1(_1755_),
    .A2(_1759_));
 sg13g2_mux4_1 _5669_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[641]),
    .A1(rf_reg[673]),
    .A2(rf_reg[705]),
    .A3(rf_reg[737]),
    .S1(raddr_a_i[1]),
    .X(_1761_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5670_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[513]),
    .A1(rf_reg[545]),
    .A2(rf_reg[577]),
    .A3(rf_reg[609]),
    .S1(raddr_a_i[1]),
    .X(_1762_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5671_ (.A0(rf_reg[449]),
    .A1(rf_reg[481]),
    .S(raddr_a_i[0]),
    .X(_1763_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5672_ (.A0(rf_reg[385]),
    .A1(rf_reg[417]),
    .S(raddr_a_i[0]),
    .X(_1764_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5673_ (.Y(_1765_),
    .B1(_1764_),
    .B2(net267),
    .A2(_1763_),
    .A1(net283),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5674_ (.A0(rf_reg[321]),
    .A1(rf_reg[353]),
    .S(raddr_a_i[0]),
    .X(_1766_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5675_ (.A0(rf_reg[257]),
    .A1(rf_reg[289]),
    .S(raddr_a_i[0]),
    .X(_1767_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5676_ (.Y(_1768_),
    .B1(_1767_),
    .B2(net253),
    .A2(_1766_),
    .A1(net242),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5677_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net235),
    .Y(_1769_),
    .A2(_1768_),
    .A1(_1765_));
 sg13g2_a221oi_1 _5678_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1769_),
    .B1(_1762_),
    .A1(net69),
    .Y(_1770_),
    .A2(_1761_));
 sg13g2_nand3_1 _5679_ (.B(_1760_),
    .C(_1770_),
    .A(_1751_),
    .Y(rdata_a_o[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5680_ (.A0(rf_reg[896]),
    .A1(rf_reg[928]),
    .S(raddr_a_i[0]),
    .X(_1771_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5681_ (.A0(rf_reg[960]),
    .A1(rf_reg[992]),
    .S(raddr_a_i[0]),
    .X(_1772_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5682_ (.Y(_1773_),
    .B1(_1772_),
    .B2(net284),
    .A2(_1771_),
    .A1(net268),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5683_ (.A0(rf_reg[768]),
    .A1(rf_reg[800]),
    .S(raddr_a_i[0]),
    .X(_1774_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5684_ (.A0(rf_reg[832]),
    .A1(rf_reg[864]),
    .S(raddr_a_i[0]),
    .X(_1775_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5685_ (.Y(_1776_),
    .B1(_1775_),
    .B2(net242),
    .A2(_1774_),
    .A1(net253),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5686_ (.A2(_1776_),
    .A1(_1773_),
    .B1(net309),
    .X(_1777_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5687_ (.A0(rf_reg[32]),
    .A1(rf_reg[96]),
    .S(raddr_a_i[1]),
    .X(_1778_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5688_ (.Y(_1779_),
    .A(raddr_a_i[0]),
    .B(_1778_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5689_ (.B(rf_reg[64]),
    .C(raddr_a_i[1]),
    .Y(_1780_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5690_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1779_),
    .A2(_1780_),
    .Y(_1781_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5691_ (.A0(rf_reg[128]),
    .A1(rf_reg[160]),
    .S(raddr_a_i[0]),
    .X(_1782_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5692_ (.A0(rf_reg[192]),
    .A1(rf_reg[224]),
    .S(raddr_a_i[0]),
    .X(_1783_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5693_ (.Y(_1784_),
    .B1(_1783_),
    .B2(net289),
    .A2(_1782_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5694_ (.VDD(VDD),
    .Y(_1785_),
    .A(_1784_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5695_ (.B1(net314),
    .VDD(VDD),
    .Y(_1786_),
    .VSS(VSS),
    .A1(_1781_),
    .A2(_1785_));
 sg13g2_mux4_1 _5696_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[640]),
    .A1(rf_reg[672]),
    .A2(rf_reg[704]),
    .A3(rf_reg[736]),
    .S1(raddr_a_i[1]),
    .X(_1787_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5697_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[512]),
    .A1(rf_reg[544]),
    .A2(rf_reg[576]),
    .A3(rf_reg[608]),
    .S1(raddr_a_i[1]),
    .X(_1788_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5698_ (.A0(rf_reg[448]),
    .A1(rf_reg[480]),
    .S(raddr_a_i[0]),
    .X(_1789_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5699_ (.A0(rf_reg[384]),
    .A1(rf_reg[416]),
    .S(raddr_a_i[0]),
    .X(_1790_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5700_ (.Y(_1791_),
    .B1(_1790_),
    .B2(net267),
    .A2(_1789_),
    .A1(net283),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5701_ (.A0(rf_reg[320]),
    .A1(rf_reg[352]),
    .S(raddr_a_i[0]),
    .X(_1792_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5702_ (.A0(rf_reg[256]),
    .A1(rf_reg[288]),
    .S(raddr_a_i[0]),
    .X(_1793_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5703_ (.Y(_1794_),
    .B1(_1793_),
    .B2(net253),
    .A2(_1792_),
    .A1(net242),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5704_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net235),
    .Y(_1795_),
    .A2(_1794_),
    .A1(_1791_));
 sg13g2_a221oi_1 _5705_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net230),
    .C1(_1795_),
    .B1(_1788_),
    .A1(net69),
    .Y(_1796_),
    .A2(_1787_));
 sg13g2_nand3_1 _5706_ (.B(_1786_),
    .C(_1796_),
    .A(_1777_),
    .Y(rdata_a_o[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5707_ (.A0(rf_reg[923]),
    .A1(rf_reg[955]),
    .S(raddr_a_i[0]),
    .X(_1797_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5708_ (.A0(rf_reg[987]),
    .A1(rf_reg[1019]),
    .S(raddr_a_i[0]),
    .X(_1798_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5709_ (.Y(_1799_),
    .B1(_1798_),
    .B2(net284),
    .A2(_1797_),
    .A1(net268),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5710_ (.A0(rf_reg[795]),
    .A1(rf_reg[827]),
    .S(raddr_a_i[0]),
    .X(_1800_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5711_ (.A0(rf_reg[859]),
    .A1(rf_reg[891]),
    .S(raddr_a_i[0]),
    .X(_1801_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5712_ (.Y(_1802_),
    .B1(_1801_),
    .B2(net245),
    .A2(_1800_),
    .A1(net254),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5713_ (.A2(_1802_),
    .A1(_1799_),
    .B1(net310),
    .X(_1803_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5714_ (.A0(rf_reg[59]),
    .A1(rf_reg[123]),
    .S(raddr_a_i[1]),
    .X(_1804_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5715_ (.Y(_1805_),
    .A(raddr_a_i[0]),
    .B(_1804_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5716_ (.B(rf_reg[91]),
    .C(raddr_a_i[1]),
    .Y(_1806_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5717_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1805_),
    .A2(_1806_),
    .Y(_1807_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5718_ (.A0(rf_reg[155]),
    .A1(rf_reg[187]),
    .S(raddr_a_i[0]),
    .X(_1808_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5719_ (.A0(rf_reg[219]),
    .A1(rf_reg[251]),
    .S(raddr_a_i[0]),
    .X(_1809_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5720_ (.Y(_1810_),
    .B1(_1809_),
    .B2(net289),
    .A2(_1808_),
    .A1(net273),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5721_ (.VDD(VDD),
    .Y(_1811_),
    .A(_1810_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5722_ (.B1(net313),
    .VDD(VDD),
    .Y(_1812_),
    .VSS(VSS),
    .A1(_1807_),
    .A2(_1811_));
 sg13g2_mux4_1 _5723_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[667]),
    .A1(rf_reg[699]),
    .A2(rf_reg[731]),
    .A3(rf_reg[763]),
    .S1(raddr_a_i[1]),
    .X(_1813_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5724_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[539]),
    .A1(rf_reg[571]),
    .A2(rf_reg[603]),
    .A3(rf_reg[635]),
    .S1(raddr_a_i[1]),
    .X(_1814_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5725_ (.A0(rf_reg[475]),
    .A1(rf_reg[507]),
    .S(raddr_a_i[0]),
    .X(_1815_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5726_ (.A0(rf_reg[411]),
    .A1(rf_reg[443]),
    .S(raddr_a_i[0]),
    .X(_1816_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5727_ (.Y(_1817_),
    .B1(_1816_),
    .B2(net270),
    .A2(_1815_),
    .A1(net286),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5728_ (.A0(rf_reg[347]),
    .A1(rf_reg[379]),
    .S(raddr_a_i[0]),
    .X(_1818_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5729_ (.A0(rf_reg[283]),
    .A1(rf_reg[315]),
    .S(raddr_a_i[0]),
    .X(_1819_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5730_ (.Y(_1820_),
    .B1(_1819_),
    .B2(net256),
    .A2(_1818_),
    .A1(net245),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5731_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1817_),
    .A2(_1820_),
    .Y(_1821_),
    .B1(net236));
 sg13g2_a221oi_1 _5732_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1821_),
    .B1(_1814_),
    .A1(net68),
    .Y(_1822_),
    .A2(_1813_));
 sg13g2_nand3_1 _5733_ (.B(_1812_),
    .C(_1822_),
    .A(_1803_),
    .Y(rdata_a_o[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5734_ (.A0(rf_reg[922]),
    .A1(rf_reg[954]),
    .S(raddr_a_i[0]),
    .X(_1823_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5735_ (.A0(rf_reg[986]),
    .A1(rf_reg[1018]),
    .S(raddr_a_i[0]),
    .X(_1824_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5736_ (.Y(_1825_),
    .B1(_1824_),
    .B2(net275),
    .A2(_1823_),
    .A1(net259),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5737_ (.A0(rf_reg[794]),
    .A1(rf_reg[826]),
    .S(raddr_a_i[0]),
    .X(_1826_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5738_ (.A0(rf_reg[858]),
    .A1(rf_reg[890]),
    .S(raddr_a_i[0]),
    .X(_1827_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5739_ (.Y(_1828_),
    .B1(_1827_),
    .B2(net238),
    .A2(_1826_),
    .A1(net249),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5740_ (.A2(_1828_),
    .A1(_1825_),
    .B1(net306),
    .X(_1829_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5741_ (.A0(rf_reg[58]),
    .A1(rf_reg[122]),
    .S(raddr_a_i[1]),
    .X(_1830_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5742_ (.Y(_1831_),
    .A(raddr_a_i[0]),
    .B(_1830_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5743_ (.B(rf_reg[90]),
    .C(raddr_a_i[1]),
    .Y(_1832_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5744_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1831_),
    .A2(_1832_),
    .Y(_1833_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5745_ (.A0(rf_reg[154]),
    .A1(rf_reg[186]),
    .S(raddr_a_i[0]),
    .X(_1834_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5746_ (.A0(rf_reg[218]),
    .A1(rf_reg[250]),
    .S(raddr_a_i[0]),
    .X(_1835_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5747_ (.Y(_1836_),
    .B1(_1835_),
    .B2(net280),
    .A2(_1834_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5748_ (.VDD(VDD),
    .Y(_1837_),
    .A(_1836_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5749_ (.B1(net312),
    .VDD(VDD),
    .Y(_1838_),
    .VSS(VSS),
    .A1(_1833_),
    .A2(_1837_));
 sg13g2_mux4_1 _5750_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[666]),
    .A1(rf_reg[698]),
    .A2(rf_reg[730]),
    .A3(rf_reg[762]),
    .S1(raddr_a_i[1]),
    .X(_1839_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5751_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[538]),
    .A1(rf_reg[570]),
    .A2(rf_reg[602]),
    .A3(rf_reg[634]),
    .S1(raddr_a_i[1]),
    .X(_1840_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5752_ (.A0(rf_reg[474]),
    .A1(rf_reg[506]),
    .S(raddr_a_i[0]),
    .X(_1841_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5753_ (.A0(rf_reg[410]),
    .A1(rf_reg[442]),
    .S(raddr_a_i[0]),
    .X(_1842_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5754_ (.Y(_1843_),
    .B1(_1842_),
    .B2(net259),
    .A2(_1841_),
    .A1(net275),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5755_ (.A0(rf_reg[346]),
    .A1(rf_reg[378]),
    .S(raddr_a_i[0]),
    .X(_1844_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5756_ (.A0(rf_reg[282]),
    .A1(rf_reg[314]),
    .S(raddr_a_i[0]),
    .X(_1845_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5757_ (.Y(_1846_),
    .B1(_1845_),
    .B2(net249),
    .A2(_1844_),
    .A1(net238),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5758_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net232),
    .Y(_1847_),
    .A2(_1846_),
    .A1(_1843_));
 sg13g2_a221oi_1 _5759_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1847_),
    .B1(_1840_),
    .A1(net66),
    .Y(_1848_),
    .A2(_1839_));
 sg13g2_nand3_1 _5760_ (.B(_1838_),
    .C(_1848_),
    .A(_1829_),
    .Y(rdata_a_o[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5761_ (.A0(rf_reg[921]),
    .A1(rf_reg[953]),
    .S(raddr_a_i[0]),
    .X(_1849_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5762_ (.A0(rf_reg[985]),
    .A1(rf_reg[1017]),
    .S(raddr_a_i[0]),
    .X(_1850_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5763_ (.Y(_1851_),
    .B1(_1850_),
    .B2(net278),
    .A2(_1849_),
    .A1(net263),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5764_ (.A0(rf_reg[793]),
    .A1(rf_reg[825]),
    .S(raddr_a_i[0]),
    .X(_1852_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5765_ (.A0(rf_reg[857]),
    .A1(rf_reg[889]),
    .S(raddr_a_i[0]),
    .X(_1853_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5766_ (.Y(_1854_),
    .B1(_1853_),
    .B2(net240),
    .A2(_1852_),
    .A1(net251),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5767_ (.A2(_1854_),
    .A1(_1851_),
    .B1(net310),
    .X(_1855_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5768_ (.A0(rf_reg[57]),
    .A1(rf_reg[121]),
    .S(raddr_a_i[1]),
    .X(_1856_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5769_ (.Y(_1857_),
    .A(raddr_a_i[0]),
    .B(_1856_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5770_ (.B(rf_reg[89]),
    .C(raddr_a_i[1]),
    .Y(_1858_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5771_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1857_),
    .A2(_1858_),
    .Y(_1859_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5772_ (.A0(rf_reg[153]),
    .A1(rf_reg[185]),
    .S(raddr_a_i[0]),
    .X(_1860_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5773_ (.A0(rf_reg[217]),
    .A1(rf_reg[249]),
    .S(raddr_a_i[0]),
    .X(_1861_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5774_ (.Y(_1862_),
    .B1(_1861_),
    .B2(net281),
    .A2(_1860_),
    .A1(net265),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5775_ (.VDD(VDD),
    .Y(_1863_),
    .A(_1862_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5776_ (.B1(net315),
    .VDD(VDD),
    .Y(_1864_),
    .VSS(VSS),
    .A1(_1859_),
    .A2(_1863_));
 sg13g2_mux4_1 _5777_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[665]),
    .A1(rf_reg[697]),
    .A2(rf_reg[729]),
    .A3(rf_reg[761]),
    .S1(raddr_a_i[1]),
    .X(_1865_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5778_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[537]),
    .A1(rf_reg[569]),
    .A2(rf_reg[601]),
    .A3(rf_reg[633]),
    .S1(raddr_a_i[1]),
    .X(_1866_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5779_ (.A0(rf_reg[473]),
    .A1(rf_reg[505]),
    .S(raddr_a_i[0]),
    .X(_1867_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5780_ (.A0(rf_reg[409]),
    .A1(rf_reg[441]),
    .S(raddr_a_i[0]),
    .X(_1868_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5781_ (.Y(_1869_),
    .B1(_1868_),
    .B2(net261),
    .A2(_1867_),
    .A1(net277),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5782_ (.A0(rf_reg[345]),
    .A1(rf_reg[377]),
    .S(raddr_a_i[0]),
    .X(_1870_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5783_ (.A0(rf_reg[281]),
    .A1(rf_reg[313]),
    .S(raddr_a_i[0]),
    .X(_1871_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5784_ (.Y(_1872_),
    .B1(_1871_),
    .B2(net250),
    .A2(_1870_),
    .A1(net239),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5785_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net233),
    .Y(_1873_),
    .A2(_1872_),
    .A1(_1869_));
 sg13g2_a221oi_1 _5786_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net231),
    .C1(_1873_),
    .B1(_1866_),
    .A1(net70),
    .Y(_1874_),
    .A2(_1865_));
 sg13g2_nand3_1 _5787_ (.B(_1864_),
    .C(_1874_),
    .A(_1855_),
    .Y(rdata_a_o[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5788_ (.A0(rf_reg[920]),
    .A1(rf_reg[952]),
    .S(raddr_a_i[0]),
    .X(_1875_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5789_ (.A0(rf_reg[984]),
    .A1(rf_reg[1016]),
    .S(raddr_a_i[0]),
    .X(_1876_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5790_ (.Y(_1877_),
    .B1(_1876_),
    .B2(net286),
    .A2(_1875_),
    .A1(net270),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5791_ (.A0(rf_reg[792]),
    .A1(rf_reg[824]),
    .S(raddr_a_i[0]),
    .X(_1878_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5792_ (.A0(rf_reg[856]),
    .A1(rf_reg[888]),
    .S(raddr_a_i[0]),
    .X(_1879_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5793_ (.Y(_1880_),
    .B1(_1879_),
    .B2(net245),
    .A2(_1878_),
    .A1(net256),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_2 _5794_ (.A2(_1880_),
    .A1(_1877_),
    .B1(net308),
    .X(_1881_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5795_ (.A0(rf_reg[56]),
    .A1(rf_reg[120]),
    .S(raddr_a_i[1]),
    .X(_1882_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5796_ (.Y(_1883_),
    .A(raddr_a_i[0]),
    .B(_1882_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5797_ (.B(rf_reg[88]),
    .C(raddr_a_i[1]),
    .Y(_1884_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5798_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1883_),
    .A2(_1884_),
    .Y(_1885_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5799_ (.A0(rf_reg[152]),
    .A1(rf_reg[184]),
    .S(raddr_a_i[0]),
    .X(_1886_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5800_ (.A0(rf_reg[216]),
    .A1(rf_reg[248]),
    .S(raddr_a_i[0]),
    .X(_1887_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5801_ (.Y(_1888_),
    .B1(_1887_),
    .B2(net288),
    .A2(_1886_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5802_ (.VDD(VDD),
    .Y(_1889_),
    .A(_1888_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5803_ (.B1(net313),
    .VDD(VDD),
    .Y(_1890_),
    .VSS(VSS),
    .A1(_1885_),
    .A2(_1889_));
 sg13g2_mux4_1 _5804_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[664]),
    .A1(rf_reg[696]),
    .A2(rf_reg[728]),
    .A3(rf_reg[760]),
    .S1(raddr_a_i[1]),
    .X(_1891_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5805_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[536]),
    .A1(rf_reg[568]),
    .A2(rf_reg[600]),
    .A3(rf_reg[632]),
    .S1(raddr_a_i[1]),
    .X(_1892_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5806_ (.A0(rf_reg[472]),
    .A1(rf_reg[504]),
    .S(raddr_a_i[0]),
    .X(_1893_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5807_ (.A0(rf_reg[408]),
    .A1(rf_reg[440]),
    .S(raddr_a_i[0]),
    .X(_1894_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5808_ (.Y(_1895_),
    .B1(_1894_),
    .B2(net269),
    .A2(_1893_),
    .A1(net285),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5809_ (.A0(rf_reg[344]),
    .A1(rf_reg[376]),
    .S(raddr_a_i[0]),
    .X(_1896_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5810_ (.A0(rf_reg[280]),
    .A1(rf_reg[312]),
    .S(raddr_a_i[0]),
    .X(_1897_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5811_ (.Y(_1898_),
    .B1(_1897_),
    .B2(net255),
    .A2(_1896_),
    .A1(net244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5812_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net234),
    .Y(_1899_),
    .A2(_1898_),
    .A1(_1895_));
 sg13g2_a221oi_1 _5813_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1899_),
    .B1(_1892_),
    .A1(net68),
    .Y(_1900_),
    .A2(_1891_));
 sg13g2_nand3_1 _5814_ (.B(_1890_),
    .C(_1900_),
    .A(_1881_),
    .Y(rdata_a_o[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5815_ (.A0(rf_reg[919]),
    .A1(rf_reg[951]),
    .S(raddr_a_i[0]),
    .X(_1901_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5816_ (.A0(rf_reg[983]),
    .A1(rf_reg[1015]),
    .S(raddr_a_i[0]),
    .X(_1902_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5817_ (.Y(_1903_),
    .B1(_1902_),
    .B2(net286),
    .A2(_1901_),
    .A1(net270),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5818_ (.A0(rf_reg[791]),
    .A1(rf_reg[823]),
    .S(raddr_a_i[0]),
    .X(_1904_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5819_ (.A0(rf_reg[855]),
    .A1(rf_reg[887]),
    .S(raddr_a_i[0]),
    .X(_1905_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5820_ (.Y(_1906_),
    .B1(_1905_),
    .B2(net245),
    .A2(_1904_),
    .A1(net256),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5821_ (.A2(_1906_),
    .A1(_1903_),
    .B1(net308),
    .X(_1907_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5822_ (.A0(rf_reg[55]),
    .A1(rf_reg[119]),
    .S(raddr_a_i[1]),
    .X(_1908_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5823_ (.Y(_1909_),
    .A(raddr_a_i[0]),
    .B(_1908_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5824_ (.B(rf_reg[87]),
    .C(raddr_a_i[1]),
    .Y(_1910_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5825_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1909_),
    .A2(_1910_),
    .Y(_1911_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5826_ (.A0(rf_reg[151]),
    .A1(rf_reg[183]),
    .S(raddr_a_i[0]),
    .X(_1912_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5827_ (.A0(rf_reg[215]),
    .A1(rf_reg[247]),
    .S(raddr_a_i[0]),
    .X(_1913_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5828_ (.Y(_1914_),
    .B1(_1913_),
    .B2(net288),
    .A2(_1912_),
    .A1(net272),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5829_ (.VDD(VDD),
    .Y(_1915_),
    .A(_1914_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5830_ (.B1(net313),
    .VDD(VDD),
    .Y(_1916_),
    .VSS(VSS),
    .A1(_1911_),
    .A2(_1915_));
 sg13g2_mux4_1 _5831_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[663]),
    .A1(rf_reg[695]),
    .A2(rf_reg[727]),
    .A3(rf_reg[759]),
    .S1(raddr_a_i[1]),
    .X(_1917_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5832_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[535]),
    .A1(rf_reg[567]),
    .A2(rf_reg[599]),
    .A3(rf_reg[631]),
    .S1(raddr_a_i[1]),
    .X(_1918_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5833_ (.A0(rf_reg[471]),
    .A1(rf_reg[503]),
    .S(raddr_a_i[0]),
    .X(_1919_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5834_ (.A0(rf_reg[407]),
    .A1(rf_reg[439]),
    .S(raddr_a_i[0]),
    .X(_1920_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5835_ (.Y(_1921_),
    .B1(_1920_),
    .B2(net269),
    .A2(_1919_),
    .A1(net285),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5836_ (.A0(rf_reg[343]),
    .A1(rf_reg[375]),
    .S(raddr_a_i[0]),
    .X(_1922_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5837_ (.A0(rf_reg[279]),
    .A1(rf_reg[311]),
    .S(raddr_a_i[0]),
    .X(_1923_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5838_ (.Y(_1924_),
    .B1(_1923_),
    .B2(net255),
    .A2(_1922_),
    .A1(net244),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _5839_ (.VSS(VSS),
    .VDD(VDD),
    .B1(net234),
    .Y(_1925_),
    .A2(_1924_),
    .A1(_1921_));
 sg13g2_a221oi_1 _5840_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net229),
    .C1(_1925_),
    .B1(_1918_),
    .A1(net68),
    .Y(_1926_),
    .A2(_1917_));
 sg13g2_nand3_1 _5841_ (.B(_1916_),
    .C(_1926_),
    .A(_1907_),
    .Y(rdata_a_o[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5842_ (.A0(rf_reg[918]),
    .A1(rf_reg[950]),
    .S(raddr_a_i[0]),
    .X(_1927_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5843_ (.A0(rf_reg[982]),
    .A1(rf_reg[1014]),
    .S(raddr_a_i[0]),
    .X(_1928_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5844_ (.Y(_1929_),
    .B1(_1928_),
    .B2(net276),
    .A2(_1927_),
    .A1(net260),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5845_ (.A0(rf_reg[790]),
    .A1(rf_reg[822]),
    .S(raddr_a_i[0]),
    .X(_1930_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5846_ (.A0(rf_reg[854]),
    .A1(rf_reg[886]),
    .S(raddr_a_i[0]),
    .X(_1931_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5847_ (.Y(_1932_),
    .B1(_1931_),
    .B2(net237),
    .A2(_1930_),
    .A1(net248),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _5848_ (.A2(_1932_),
    .A1(_1929_),
    .B1(net306),
    .X(_1933_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5849_ (.A0(rf_reg[54]),
    .A1(rf_reg[118]),
    .S(raddr_a_i[1]),
    .X(_1934_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5850_ (.Y(_1935_),
    .A(raddr_a_i[0]),
    .B(_1934_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _5851_ (.B(rf_reg[86]),
    .C(raddr_a_i[1]),
    .Y(_1936_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(raddr_a_i[0]));
 sg13g2_a21oi_1 _5852_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1935_),
    .A2(_1936_),
    .Y(_1937_),
    .B1(raddr_a_i[2]));
 sg13g2_mux2_1 _5853_ (.A0(rf_reg[150]),
    .A1(rf_reg[182]),
    .S(raddr_a_i[0]),
    .X(_1938_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5854_ (.A0(rf_reg[214]),
    .A1(rf_reg[246]),
    .S(raddr_a_i[0]),
    .X(_1939_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5855_ (.Y(_1940_),
    .B1(_1939_),
    .B2(net280),
    .A2(_1938_),
    .A1(net264),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5856_ (.VDD(VDD),
    .Y(_1941_),
    .A(_1940_),
    .VSS(VSS));
 sg13g2_o21ai_1 _5857_ (.B1(net311),
    .VDD(VDD),
    .Y(_1942_),
    .VSS(VSS),
    .A1(_1937_),
    .A2(_1941_));
 sg13g2_mux4_1 _5858_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[662]),
    .A1(rf_reg[694]),
    .A2(rf_reg[726]),
    .A3(rf_reg[758]),
    .S1(raddr_a_i[1]),
    .X(_1943_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5859_ (.S0(raddr_a_i[0]),
    .A0(rf_reg[534]),
    .A1(rf_reg[566]),
    .A2(rf_reg[598]),
    .A3(rf_reg[630]),
    .S1(raddr_a_i[1]),
    .X(_1944_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5860_ (.A0(rf_reg[470]),
    .A1(rf_reg[502]),
    .S(raddr_a_i[0]),
    .X(_1945_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5861_ (.A0(rf_reg[406]),
    .A1(rf_reg[438]),
    .S(raddr_a_i[0]),
    .X(_1946_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5862_ (.Y(_1947_),
    .B1(_1946_),
    .B2(net260),
    .A2(_1945_),
    .A1(net276),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5863_ (.A0(rf_reg[342]),
    .A1(rf_reg[374]),
    .S(raddr_a_i[0]),
    .X(_1948_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5864_ (.A0(rf_reg[278]),
    .A1(rf_reg[310]),
    .S(raddr_a_i[0]),
    .X(_1949_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5865_ (.Y(_1950_),
    .B1(_1949_),
    .B2(net248),
    .A2(_1948_),
    .A1(net237),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5866_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1947_),
    .A2(_1950_),
    .Y(_1951_),
    .B1(net232));
 sg13g2_a221oi_1 _5867_ (.VSS(VSS),
    .VDD(VDD),
    .B2(net227),
    .C1(_1951_),
    .B1(_1944_),
    .A1(net66),
    .Y(_1952_),
    .A2(_1943_));
 sg13g2_nand3_1 _5868_ (.B(_1942_),
    .C(_1952_),
    .A(_1933_),
    .Y(rdata_a_o[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5869_ (.VDD(VDD),
    .Y(_1953_),
    .A(raddr_b_i[4]),
    .VSS(VSS));
 sg13g2_nor3_1 _5870_ (.A(_1953_),
    .B(raddr_b_i[3]),
    .C(raddr_b_i[2]),
    .Y(_1954_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout231 (.A(_1052_),
    .X(net231),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(net231),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(net230),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net231),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout227 (.A(net228),
    .X(net227),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout226 (.A(_1954_),
    .X(net226),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(net226),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5878_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[543]),
    .A1(rf_reg[575]),
    .A2(rf_reg[607]),
    .A3(rf_reg[639]),
    .S1(raddr_b_i[1]),
    .X(_1962_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _5879_ (.VDD(VDD),
    .Y(_1963_),
    .A(raddr_b_i[2]),
    .VSS(VSS));
 sg13g2_nor3_1 _5880_ (.A(_1953_),
    .B(raddr_b_i[3]),
    .C(_1963_),
    .Y(_1964_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(net226),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout221 (.A(_1964_),
    .X(net221),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5885_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[671]),
    .A1(rf_reg[703]),
    .A2(rf_reg[735]),
    .A3(rf_reg[767]),
    .S1(raddr_b_i[1]),
    .X(_1969_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5886_ (.Y(_1970_),
    .B1(net218),
    .B2(_1969_),
    .A2(_1962_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _5887_ (.VSS(VSS),
    .VDD(VDD),
    .X(_1971_),
    .B(raddr_b_i[3]),
    .A(raddr_b_i[4]));
 sg13g2_nor2_1 _5888_ (.A(raddr_b_i[2]),
    .B(net304),
    .Y(_1972_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(net221),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(net220),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(net221),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(net218),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout216 (.A(_1972_),
    .X(net216),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(net216),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5895_ (.Y(_1979_),
    .A(rf_reg[63]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(net215),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(net216),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5898_ (.A0(rf_reg[95]),
    .A1(rf_reg[127]),
    .S(raddr_b_i[0]),
    .X(_1982_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5899_ (.Y(_1983_),
    .A(raddr_b_i[1]),
    .B(_1982_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _5900_ (.B1(_1983_),
    .VDD(VDD),
    .Y(_1984_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_1979_));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(net213),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 _5902_ (.A(raddr_b_i[1]),
    .B_N(raddr_b_i[2]),
    .Y(_1986_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(_1986_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(net211),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5905_ (.A0(rf_reg[159]),
    .A1(rf_reg[191]),
    .S(raddr_b_i[0]),
    .X(_1989_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout208 (.A(net211),
    .X(net208),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5908_ (.A0(rf_reg[223]),
    .A1(rf_reg[255]),
    .S(raddr_b_i[0]),
    .X(_1992_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _5909_ (.A(raddr_b_i[1]),
    .B(raddr_b_i[2]),
    .X(_1993_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net208),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net207),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(net208),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5913_ (.Y(_1997_),
    .B1(_1992_),
    .B2(net187),
    .A2(_1989_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _5914_ (.A(net302),
    .B(_1997_),
    .Y(_1998_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5915_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_1984_),
    .Y(_1999_),
    .B1(_1998_));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net205),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(_1986_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5918_ (.A0(rf_reg[479]),
    .A1(rf_reg[511]),
    .S(raddr_b_i[0]),
    .X(_2002_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout201 (.A(_1986_),
    .X(net201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5921_ (.A0(rf_reg[351]),
    .A1(rf_reg[383]),
    .S(raddr_b_i[0]),
    .X(_2005_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 _5922_ (.A(raddr_b_i[2]),
    .B_N(raddr_b_i[1]),
    .Y(_2006_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(net201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5925_ (.Y(_2009_),
    .B1(_2005_),
    .B2(net175),
    .A2(_2002_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5926_ (.A0(rf_reg[415]),
    .A1(rf_reg[447]),
    .S(raddr_b_i[0]),
    .X(_2010_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(net201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(net201),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5929_ (.A0(rf_reg[287]),
    .A1(rf_reg[319]),
    .S(raddr_b_i[0]),
    .X(_2013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _5930_ (.A(raddr_b_i[1]),
    .B(raddr_b_i[2]),
    .Y(_2014_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(_1993_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(net196),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5933_ (.Y(_2017_),
    .B1(_2013_),
    .B2(net163),
    .A2(net199),
    .A1(_2010_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5934_ (.Y(_2018_),
    .A(_2009_),
    .B(_2017_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _5935_ (.A(raddr_b_i[4]),
    .B_N(raddr_b_i[3]),
    .Y(_2019_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(net196),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5937_ (.A0(rf_reg[927]),
    .A1(rf_reg[959]),
    .S(raddr_b_i[0]),
    .X(_2021_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(net196),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5939_ (.A0(rf_reg[799]),
    .A1(rf_reg[831]),
    .S(raddr_b_i[0]),
    .X(_2023_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(net193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5941_ (.Y(_2025_),
    .B1(_2023_),
    .B2(net163),
    .A2(_2021_),
    .A1(net199),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(net193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout190 (.A(net196),
    .X(net190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5944_ (.A0(rf_reg[863]),
    .A1(rf_reg[895]),
    .S(raddr_b_i[0]),
    .X(_2028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(net196),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5946_ (.A0(rf_reg[991]),
    .A1(rf_reg[1023]),
    .S(raddr_b_i[0]),
    .X(_2030_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(_1993_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5948_ (.Y(_2032_),
    .B1(_2030_),
    .B2(net184),
    .A2(_2028_),
    .A1(net175),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5949_ (.Y(_2033_),
    .A(_2025_),
    .B(_2032_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _5950_ (.A(raddr_b_i[4]),
    .B(raddr_b_i[3]),
    .X(_2034_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(net188),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(net187),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5953_ (.Y(_2037_),
    .B1(_2033_),
    .B2(net292),
    .A2(net297),
    .A1(_2018_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _5954_ (.B(_1999_),
    .C(_2037_),
    .A(_1970_),
    .Y(rdata_b_o[31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5955_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[542]),
    .A1(rf_reg[574]),
    .A2(rf_reg[606]),
    .A3(rf_reg[638]),
    .S1(raddr_b_i[1]),
    .X(_2038_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5956_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[670]),
    .A1(rf_reg[702]),
    .A2(rf_reg[734]),
    .A3(rf_reg[766]),
    .S1(raddr_b_i[1]),
    .X(_2039_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(net188),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5958_ (.Y(_2041_),
    .B1(_2039_),
    .B2(net218),
    .A2(_2038_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5959_ (.Y(_2042_),
    .A(rf_reg[62]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5960_ (.A0(rf_reg[94]),
    .A1(rf_reg[126]),
    .S(raddr_b_i[0]),
    .X(_2043_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5961_ (.Y(_2044_),
    .A(raddr_b_i[1]),
    .B(_2043_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _5962_ (.B1(_2044_),
    .VDD(VDD),
    .Y(_2045_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2042_));
 sg13g2_mux2_1 _5963_ (.A0(rf_reg[158]),
    .A1(rf_reg[190]),
    .S(raddr_b_i[0]),
    .X(_2046_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5964_ (.A0(rf_reg[222]),
    .A1(rf_reg[254]),
    .S(raddr_b_i[0]),
    .X(_2047_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5965_ (.Y(_2048_),
    .B1(_2047_),
    .B2(net187),
    .A2(_2046_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _5966_ (.A(net302),
    .B(_2048_),
    .Y(_2049_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5967_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_2045_),
    .Y(_2050_),
    .B1(_2049_));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5969_ (.A0(rf_reg[478]),
    .A1(rf_reg[510]),
    .S(raddr_b_i[0]),
    .X(_2052_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(net188),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5971_ (.A0(rf_reg[350]),
    .A1(rf_reg[382]),
    .S(raddr_b_i[0]),
    .X(_2054_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5972_ (.Y(_2055_),
    .B1(_2054_),
    .B2(net176),
    .A2(_2052_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5973_ (.A0(rf_reg[414]),
    .A1(rf_reg[446]),
    .S(raddr_b_i[0]),
    .X(_2056_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5974_ (.A0(rf_reg[286]),
    .A1(rf_reg[318]),
    .S(raddr_b_i[0]),
    .X(_2057_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5975_ (.Y(_2058_),
    .B1(_2057_),
    .B2(net164),
    .A2(_2056_),
    .A1(net200),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5976_ (.Y(_2059_),
    .A(_2055_),
    .B(_2058_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5977_ (.A0(rf_reg[990]),
    .A1(rf_reg[1022]),
    .S(raddr_b_i[0]),
    .X(_2060_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5978_ (.A0(rf_reg[798]),
    .A1(rf_reg[830]),
    .S(raddr_b_i[0]),
    .X(_2061_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5979_ (.Y(_2062_),
    .B1(_2061_),
    .B2(net164),
    .A2(_2060_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5980_ (.A0(rf_reg[862]),
    .A1(rf_reg[894]),
    .S(raddr_b_i[0]),
    .X(_2063_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5981_ (.A0(rf_reg[926]),
    .A1(rf_reg[958]),
    .S(raddr_b_i[0]),
    .X(_2064_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net188),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_2006_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5984_ (.Y(_2067_),
    .B1(_2064_),
    .B2(net200),
    .A2(_2063_),
    .A1(net176),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5985_ (.Y(_2068_),
    .A(_2062_),
    .B(_2067_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5986_ (.Y(_2069_),
    .B1(_2068_),
    .B2(net292),
    .A2(_2059_),
    .A1(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _5987_ (.B(_2050_),
    .C(_2069_),
    .A(_2041_),
    .Y(rdata_b_o[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5988_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[533]),
    .A1(rf_reg[565]),
    .A2(rf_reg[597]),
    .A3(rf_reg[629]),
    .S1(raddr_b_i[1]),
    .X(_2070_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _5989_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[661]),
    .A1(rf_reg[693]),
    .A2(rf_reg[725]),
    .A3(rf_reg[757]),
    .S1(raddr_b_i[1]),
    .X(_2071_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5990_ (.Y(_2072_),
    .B1(_2071_),
    .B2(net217),
    .A2(_2070_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5991_ (.Y(_2073_),
    .A(rf_reg[53]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5992_ (.A0(rf_reg[85]),
    .A1(rf_reg[117]),
    .S(raddr_b_i[0]),
    .X(_2074_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _5993_ (.Y(_2075_),
    .A(raddr_b_i[1]),
    .B(_2074_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _5994_ (.B1(_2075_),
    .VDD(VDD),
    .Y(_2076_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2073_));
 sg13g2_mux2_1 _5995_ (.A0(rf_reg[149]),
    .A1(rf_reg[181]),
    .S(raddr_b_i[0]),
    .X(_2077_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _5996_ (.A0(rf_reg[213]),
    .A1(rf_reg[245]),
    .S(raddr_b_i[0]),
    .X(_2078_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _5997_ (.Y(_2079_),
    .B1(_2078_),
    .B2(net186),
    .A2(_2077_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _5998_ (.A(net301),
    .B(_2079_),
    .Y(_2080_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _5999_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2076_),
    .Y(_2081_),
    .B1(_2080_));
 sg13g2_mux2_1 _6000_ (.A0(rf_reg[469]),
    .A1(rf_reg[501]),
    .S(raddr_b_i[0]),
    .X(_2082_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6001_ (.A0(rf_reg[341]),
    .A1(rf_reg[373]),
    .S(raddr_b_i[0]),
    .X(_2083_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6002_ (.Y(_2084_),
    .B1(_2083_),
    .B2(net173),
    .A2(_2082_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6003_ (.A0(rf_reg[405]),
    .A1(rf_reg[437]),
    .S(raddr_b_i[0]),
    .X(_2085_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6004_ (.A0(rf_reg[277]),
    .A1(rf_reg[309]),
    .S(raddr_b_i[0]),
    .X(_2086_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6005_ (.Y(_2087_),
    .B1(_2086_),
    .B2(net162),
    .A2(_2085_),
    .A1(net198),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6006_ (.Y(_2088_),
    .A(_2084_),
    .B(_2087_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6007_ (.A0(rf_reg[981]),
    .A1(rf_reg[1013]),
    .S(raddr_b_i[0]),
    .X(_2089_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6008_ (.A0(rf_reg[789]),
    .A1(rf_reg[821]),
    .S(raddr_b_i[0]),
    .X(_2090_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6009_ (.Y(_2091_),
    .B1(_2090_),
    .B2(net162),
    .A2(_2089_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6010_ (.A0(rf_reg[853]),
    .A1(rf_reg[885]),
    .S(raddr_b_i[0]),
    .X(_2092_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6011_ (.A0(rf_reg[917]),
    .A1(rf_reg[949]),
    .S(raddr_b_i[0]),
    .X(_2093_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6012_ (.Y(_2094_),
    .B1(_2093_),
    .B2(net198),
    .A2(_2092_),
    .A1(net173),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6013_ (.Y(_2095_),
    .A(_2091_),
    .B(_2094_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6014_ (.Y(_2096_),
    .B1(_2095_),
    .B2(net292),
    .A2(_2088_),
    .A1(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6015_ (.B(_2081_),
    .C(_2096_),
    .A(_2072_),
    .Y(rdata_b_o[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6016_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[532]),
    .A1(rf_reg[564]),
    .A2(rf_reg[596]),
    .A3(rf_reg[628]),
    .S1(raddr_b_i[1]),
    .X(_2097_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6017_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[660]),
    .A1(rf_reg[692]),
    .A2(rf_reg[724]),
    .A3(rf_reg[756]),
    .S1(raddr_b_i[1]),
    .X(_2098_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6018_ (.Y(_2099_),
    .B1(_2098_),
    .B2(net219),
    .A2(_2097_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6019_ (.Y(_2100_),
    .A(rf_reg[52]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6020_ (.A0(rf_reg[84]),
    .A1(rf_reg[116]),
    .S(raddr_b_i[0]),
    .X(_2101_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6021_ (.Y(_2102_),
    .A(raddr_b_i[1]),
    .B(_2101_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6022_ (.B1(_2102_),
    .VDD(VDD),
    .Y(_2103_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2100_));
 sg13g2_mux2_1 _6023_ (.A0(rf_reg[148]),
    .A1(rf_reg[180]),
    .S(raddr_b_i[0]),
    .X(_2104_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6024_ (.A0(rf_reg[212]),
    .A1(rf_reg[244]),
    .S(raddr_b_i[0]),
    .X(_2105_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6025_ (.Y(_2106_),
    .B1(_2105_),
    .B2(net195),
    .A2(_2104_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6026_ (.A(net303),
    .B(_2106_),
    .Y(_2107_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6027_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2103_),
    .Y(_2108_),
    .B1(_2107_));
 sg13g2_mux2_1 _6028_ (.A0(rf_reg[468]),
    .A1(rf_reg[500]),
    .S(raddr_b_i[0]),
    .X(_2109_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6029_ (.A0(rf_reg[340]),
    .A1(rf_reg[372]),
    .S(raddr_b_i[0]),
    .X(_2110_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6030_ (.Y(_2111_),
    .B1(_2110_),
    .B2(net180),
    .A2(_2109_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6031_ (.A0(rf_reg[404]),
    .A1(rf_reg[436]),
    .S(raddr_b_i[0]),
    .X(_2112_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6032_ (.A0(rf_reg[276]),
    .A1(rf_reg[308]),
    .S(raddr_b_i[0]),
    .X(_2113_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6033_ (.Y(_2114_),
    .B1(_2113_),
    .B2(net169),
    .A2(_2112_),
    .A1(net207),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6034_ (.Y(_2115_),
    .A(_2111_),
    .B(_2114_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6035_ (.A0(rf_reg[980]),
    .A1(rf_reg[1012]),
    .S(raddr_b_i[0]),
    .X(_2116_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6036_ (.A0(rf_reg[788]),
    .A1(rf_reg[820]),
    .S(raddr_b_i[0]),
    .X(_2117_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6037_ (.Y(_2118_),
    .B1(_2117_),
    .B2(net169),
    .A2(_2116_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net181),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6039_ (.A0(rf_reg[852]),
    .A1(rf_reg[884]),
    .S(raddr_b_i[0]),
    .X(_2120_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(net181),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6041_ (.A0(rf_reg[916]),
    .A1(rf_reg[948]),
    .S(raddr_b_i[0]),
    .X(_2122_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6042_ (.Y(_2123_),
    .B1(_2122_),
    .B2(net207),
    .A2(_2120_),
    .A1(net180),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6043_ (.Y(_2124_),
    .A(_2118_),
    .B(_2123_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6044_ (.Y(_2125_),
    .B1(_2124_),
    .B2(net293),
    .A2(_2115_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6045_ (.B(_2108_),
    .C(_2125_),
    .A(_2099_),
    .Y(rdata_b_o[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout178 (.A(net181),
    .X(net178),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6047_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[531]),
    .A1(rf_reg[563]),
    .A2(rf_reg[595]),
    .A3(rf_reg[627]),
    .S1(raddr_b_i[1]),
    .X(_2127_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6048_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[659]),
    .A1(rf_reg[691]),
    .A2(rf_reg[723]),
    .A3(rf_reg[755]),
    .S1(raddr_b_i[1]),
    .X(_2128_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6049_ (.Y(_2129_),
    .B1(_2128_),
    .B2(net220),
    .A2(_2127_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6050_ (.Y(_2130_),
    .A(rf_reg[51]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6051_ (.A0(rf_reg[83]),
    .A1(rf_reg[115]),
    .S(raddr_b_i[0]),
    .X(_2131_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6052_ (.Y(_2132_),
    .A(raddr_b_i[1]),
    .B(_2131_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6053_ (.B1(_2132_),
    .VDD(VDD),
    .Y(_2133_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2130_));
 sg13g2_mux2_1 _6054_ (.A0(rf_reg[147]),
    .A1(rf_reg[179]),
    .S(raddr_b_i[0]),
    .X(_2134_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(net181),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6056_ (.A0(rf_reg[211]),
    .A1(rf_reg[243]),
    .S(raddr_b_i[0]),
    .X(_2136_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6057_ (.Y(_2137_),
    .B1(_2136_),
    .B2(net194),
    .A2(_2134_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6058_ (.A(net304),
    .B(_2137_),
    .Y(_2138_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6059_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2133_),
    .Y(_2139_),
    .B1(_2138_));
 sg13g2_mux2_1 _6060_ (.A0(rf_reg[467]),
    .A1(rf_reg[499]),
    .S(raddr_b_i[0]),
    .X(_2140_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6061_ (.A0(rf_reg[339]),
    .A1(rf_reg[371]),
    .S(raddr_b_i[0]),
    .X(_2141_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6062_ (.Y(_2142_),
    .B1(_2141_),
    .B2(net178),
    .A2(_2140_),
    .A1(net190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6063_ (.A0(rf_reg[403]),
    .A1(rf_reg[435]),
    .S(raddr_b_i[0]),
    .X(_2143_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6064_ (.A0(rf_reg[275]),
    .A1(rf_reg[307]),
    .S(raddr_b_i[0]),
    .X(_2144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6065_ (.Y(_2145_),
    .B1(_2144_),
    .B2(net167),
    .A2(_2143_),
    .A1(net205),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6066_ (.Y(_2146_),
    .A(_2142_),
    .B(_2145_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6067_ (.A0(rf_reg[979]),
    .A1(rf_reg[1011]),
    .S(raddr_b_i[0]),
    .X(_2147_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6068_ (.A0(rf_reg[787]),
    .A1(rf_reg[819]),
    .S(raddr_b_i[0]),
    .X(_2148_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6069_ (.Y(_2149_),
    .B1(_2148_),
    .B2(net167),
    .A2(_2147_),
    .A1(net190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6070_ (.A0(rf_reg[851]),
    .A1(rf_reg[883]),
    .S(raddr_b_i[0]),
    .X(_2150_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6071_ (.A0(rf_reg[915]),
    .A1(rf_reg[947]),
    .S(raddr_b_i[0]),
    .X(_2151_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6072_ (.Y(_2152_),
    .B1(_2151_),
    .B2(net205),
    .A2(_2150_),
    .A1(net178),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6073_ (.Y(_2153_),
    .A(_2149_),
    .B(_2152_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6074_ (.Y(_2154_),
    .B1(_2153_),
    .B2(net294),
    .A2(_2146_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6075_ (.B(_2139_),
    .C(_2154_),
    .A(_2129_),
    .Y(rdata_b_o[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6076_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[530]),
    .A1(rf_reg[562]),
    .A2(rf_reg[594]),
    .A3(rf_reg[626]),
    .S1(raddr_b_i[1]),
    .X(_2155_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6077_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[658]),
    .A1(rf_reg[690]),
    .A2(rf_reg[722]),
    .A3(rf_reg[754]),
    .S1(raddr_b_i[1]),
    .X(_2156_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6078_ (.Y(_2157_),
    .B1(_2156_),
    .B2(net220),
    .A2(_2155_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6079_ (.Y(_2158_),
    .A(rf_reg[50]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6080_ (.A0(rf_reg[82]),
    .A1(rf_reg[114]),
    .S(raddr_b_i[0]),
    .X(_2159_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6081_ (.Y(_2160_),
    .A(raddr_b_i[1]),
    .B(_2159_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6082_ (.B1(_2160_),
    .VDD(VDD),
    .Y(_2161_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2158_));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(_2006_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6084_ (.A0(rf_reg[146]),
    .A1(rf_reg[178]),
    .S(raddr_b_i[0]),
    .X(_2163_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6085_ (.A0(rf_reg[210]),
    .A1(rf_reg[242]),
    .S(raddr_b_i[0]),
    .X(_2164_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6086_ (.Y(_2165_),
    .B1(_2164_),
    .B2(net194),
    .A2(_2163_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6087_ (.A(net304),
    .B(_2165_),
    .Y(_2166_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6088_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2161_),
    .Y(_2167_),
    .B1(_2166_));
 sg13g2_mux2_1 _6089_ (.A0(rf_reg[466]),
    .A1(rf_reg[498]),
    .S(raddr_b_i[0]),
    .X(_2168_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6090_ (.A0(rf_reg[338]),
    .A1(rf_reg[370]),
    .S(raddr_b_i[0]),
    .X(_2169_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6091_ (.Y(_2170_),
    .B1(_2169_),
    .B2(net178),
    .A2(_2168_),
    .A1(net190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net176),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6093_ (.A0(rf_reg[402]),
    .A1(rf_reg[434]),
    .S(raddr_b_i[0]),
    .X(_2172_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout174 (.A(_2006_),
    .X(net174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6095_ (.A0(rf_reg[274]),
    .A1(rf_reg[306]),
    .S(raddr_b_i[0]),
    .X(_2174_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6096_ (.Y(_2175_),
    .B1(_2174_),
    .B2(net167),
    .A2(_2172_),
    .A1(net205),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6097_ (.Y(_2176_),
    .A(_2170_),
    .B(_2175_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6098_ (.A0(rf_reg[978]),
    .A1(rf_reg[1010]),
    .S(raddr_b_i[0]),
    .X(_2177_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6099_ (.A0(rf_reg[786]),
    .A1(rf_reg[818]),
    .S(raddr_b_i[0]),
    .X(_2178_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6100_ (.Y(_2179_),
    .B1(_2178_),
    .B2(net167),
    .A2(_2177_),
    .A1(net190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6101_ (.A0(rf_reg[850]),
    .A1(rf_reg[882]),
    .S(raddr_b_i[0]),
    .X(_2180_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6102_ (.A0(rf_reg[914]),
    .A1(rf_reg[946]),
    .S(raddr_b_i[0]),
    .X(_2181_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6103_ (.Y(_2182_),
    .B1(_2181_),
    .B2(net205),
    .A2(_2180_),
    .A1(net178),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6104_ (.Y(_2183_),
    .A(_2179_),
    .B(_2182_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6105_ (.Y(_2184_),
    .B1(_2183_),
    .B2(net294),
    .A2(_2176_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6106_ (.B(_2167_),
    .C(_2184_),
    .A(_2157_),
    .Y(rdata_b_o[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6108_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[529]),
    .A1(rf_reg[561]),
    .A2(rf_reg[593]),
    .A3(rf_reg[625]),
    .S1(raddr_b_i[1]),
    .X(_2186_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6109_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[657]),
    .A1(rf_reg[689]),
    .A2(rf_reg[721]),
    .A3(rf_reg[753]),
    .S1(raddr_b_i[1]),
    .X(_2187_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6110_ (.Y(_2188_),
    .B1(_2187_),
    .B2(net217),
    .A2(_2186_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6111_ (.Y(_2189_),
    .A(rf_reg[49]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6113_ (.A0(rf_reg[81]),
    .A1(rf_reg[113]),
    .S(raddr_b_i[0]),
    .X(_2191_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6114_ (.Y(_2192_),
    .A(raddr_b_i[1]),
    .B(_2191_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6115_ (.B1(_2192_),
    .VDD(VDD),
    .Y(_2193_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2189_));
 sg13g2_mux2_1 _6116_ (.A0(rf_reg[145]),
    .A1(rf_reg[177]),
    .S(raddr_b_i[0]),
    .X(_2194_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6117_ (.A0(rf_reg[209]),
    .A1(rf_reg[241]),
    .S(raddr_b_i[0]),
    .X(_2195_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6118_ (.Y(_2196_),
    .B1(_2195_),
    .B2(net186),
    .A2(_2194_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6119_ (.A(net301),
    .B(_2196_),
    .Y(_2197_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6120_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2193_),
    .Y(_2198_),
    .B1(_2197_));
 sg13g2_buf_2 fanout171 (.A(_2014_),
    .X(net171),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6122_ (.A0(rf_reg[465]),
    .A1(rf_reg[497]),
    .S(raddr_b_i[0]),
    .X(_2200_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6123_ (.A0(rf_reg[337]),
    .A1(rf_reg[369]),
    .S(raddr_b_i[0]),
    .X(_2201_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6124_ (.Y(_2202_),
    .B1(_2201_),
    .B2(net173),
    .A2(_2200_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6126_ (.A0(rf_reg[401]),
    .A1(rf_reg[433]),
    .S(raddr_b_i[0]),
    .X(_2204_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6127_ (.A0(rf_reg[273]),
    .A1(rf_reg[305]),
    .S(raddr_b_i[0]),
    .X(_2205_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6128_ (.Y(_2206_),
    .B1(_2205_),
    .B2(net162),
    .A2(_2204_),
    .A1(net198),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6129_ (.Y(_2207_),
    .A(_2202_),
    .B(_2206_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6130_ (.A0(rf_reg[977]),
    .A1(rf_reg[1009]),
    .S(raddr_b_i[0]),
    .X(_2208_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6131_ (.A0(rf_reg[785]),
    .A1(rf_reg[817]),
    .S(raddr_b_i[0]),
    .X(_2209_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6132_ (.Y(_2210_),
    .B1(_2209_),
    .B2(net162),
    .A2(_2208_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6133_ (.A0(rf_reg[849]),
    .A1(rf_reg[881]),
    .S(raddr_b_i[0]),
    .X(_2211_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6134_ (.A0(rf_reg[913]),
    .A1(rf_reg[945]),
    .S(raddr_b_i[0]),
    .X(_2212_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6135_ (.Y(_2213_),
    .B1(_2212_),
    .B2(net198),
    .A2(_2211_),
    .A1(net173),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6136_ (.Y(_2214_),
    .A(_2210_),
    .B(_2213_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6137_ (.Y(_2215_),
    .B1(_2214_),
    .B2(net291),
    .A2(_2207_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6138_ (.B(_2198_),
    .C(_2215_),
    .A(_2188_),
    .Y(rdata_b_o[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6139_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[528]),
    .A1(rf_reg[560]),
    .A2(rf_reg[592]),
    .A3(rf_reg[624]),
    .S1(raddr_b_i[1]),
    .X(_2216_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6140_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[656]),
    .A1(rf_reg[688]),
    .A2(rf_reg[720]),
    .A3(rf_reg[752]),
    .S1(raddr_b_i[1]),
    .X(_2217_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6141_ (.Y(_2218_),
    .B1(_2217_),
    .B2(net219),
    .A2(_2216_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6142_ (.Y(_2219_),
    .A(rf_reg[48]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net171),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6144_ (.A0(rf_reg[80]),
    .A1(rf_reg[112]),
    .S(raddr_b_i[0]),
    .X(_2221_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6145_ (.Y(_2222_),
    .A(raddr_b_i[1]),
    .B(_2221_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6146_ (.B1(_2222_),
    .VDD(VDD),
    .Y(_2223_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2219_));
 sg13g2_mux2_1 _6147_ (.A0(rf_reg[144]),
    .A1(rf_reg[176]),
    .S(raddr_b_i[0]),
    .X(_2224_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6148_ (.A0(rf_reg[208]),
    .A1(rf_reg[240]),
    .S(raddr_b_i[0]),
    .X(_2225_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6149_ (.Y(_2226_),
    .B1(_2225_),
    .B2(net194),
    .A2(_2224_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6150_ (.A(net303),
    .B(_2226_),
    .Y(_2227_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6151_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2223_),
    .Y(_2228_),
    .B1(_2227_));
 sg13g2_mux2_1 _6152_ (.A0(rf_reg[464]),
    .A1(rf_reg[496]),
    .S(raddr_b_i[0]),
    .X(_2229_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6153_ (.A0(rf_reg[336]),
    .A1(rf_reg[368]),
    .S(raddr_b_i[0]),
    .X(_2230_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6154_ (.Y(_2231_),
    .B1(_2230_),
    .B2(net177),
    .A2(_2229_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6155_ (.A0(rf_reg[400]),
    .A1(rf_reg[432]),
    .S(raddr_b_i[0]),
    .X(_2232_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6156_ (.A0(rf_reg[272]),
    .A1(rf_reg[304]),
    .S(raddr_b_i[0]),
    .X(_2233_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6157_ (.Y(_2234_),
    .B1(_2233_),
    .B2(net166),
    .A2(_2232_),
    .A1(net204),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6158_ (.Y(_2235_),
    .A(_2231_),
    .B(_2234_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net170),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6160_ (.A0(rf_reg[976]),
    .A1(rf_reg[1008]),
    .S(raddr_b_i[0]),
    .X(_2237_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6161_ (.A0(rf_reg[784]),
    .A1(rf_reg[816]),
    .S(raddr_b_i[0]),
    .X(_2238_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6162_ (.Y(_2239_),
    .B1(_2238_),
    .B2(net169),
    .A2(_2237_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6163_ (.A0(rf_reg[848]),
    .A1(rf_reg[880]),
    .S(raddr_b_i[0]),
    .X(_2240_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6164_ (.A0(rf_reg[912]),
    .A1(rf_reg[944]),
    .S(raddr_b_i[0]),
    .X(_2241_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6165_ (.Y(_2242_),
    .B1(_2241_),
    .B2(net204),
    .A2(_2240_),
    .A1(net177),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6166_ (.Y(_2243_),
    .A(_2239_),
    .B(_2242_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6167_ (.Y(_2244_),
    .B1(_2243_),
    .B2(net293),
    .A2(_2235_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6168_ (.B(_2228_),
    .C(_2244_),
    .A(_2218_),
    .Y(rdata_b_o[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6169_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[527]),
    .A1(rf_reg[559]),
    .A2(rf_reg[591]),
    .A3(rf_reg[623]),
    .S1(raddr_b_i[1]),
    .X(_2245_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net171),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net167),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6172_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[655]),
    .A1(rf_reg[687]),
    .A2(rf_reg[719]),
    .A3(rf_reg[751]),
    .S1(raddr_b_i[1]),
    .X(_2248_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6173_ (.Y(_2249_),
    .B1(_2248_),
    .B2(net218),
    .A2(_2245_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6174_ (.Y(_2250_),
    .A(rf_reg[47]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6175_ (.A0(rf_reg[79]),
    .A1(rf_reg[111]),
    .S(raddr_b_i[0]),
    .X(_2251_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6176_ (.Y(_2252_),
    .A(raddr_b_i[1]),
    .B(_2251_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6177_ (.B1(_2252_),
    .VDD(VDD),
    .Y(_2253_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2250_));
 sg13g2_mux2_1 _6178_ (.A0(rf_reg[143]),
    .A1(rf_reg[175]),
    .S(raddr_b_i[0]),
    .X(_2254_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6179_ (.A0(rf_reg[207]),
    .A1(rf_reg[239]),
    .S(raddr_b_i[0]),
    .X(_2255_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6180_ (.Y(_2256_),
    .B1(_2255_),
    .B2(net187),
    .A2(_2254_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6181_ (.A(net302),
    .B(_2256_),
    .Y(_2257_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6182_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_2253_),
    .Y(_2258_),
    .B1(_2257_));
 sg13g2_mux2_1 _6183_ (.A0(rf_reg[463]),
    .A1(rf_reg[495]),
    .S(raddr_b_i[0]),
    .X(_2259_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6184_ (.A0(rf_reg[335]),
    .A1(rf_reg[367]),
    .S(raddr_b_i[0]),
    .X(_2260_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6185_ (.Y(_2261_),
    .B1(_2260_),
    .B2(net178),
    .A2(_2259_),
    .A1(net190),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6186_ (.A0(rf_reg[399]),
    .A1(rf_reg[431]),
    .S(raddr_b_i[0]),
    .X(_2262_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6187_ (.A0(rf_reg[271]),
    .A1(rf_reg[303]),
    .S(raddr_b_i[0]),
    .X(_2263_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout165 (.A(net171),
    .X(net165),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6189_ (.Y(_2265_),
    .B1(_2263_),
    .B2(net167),
    .A2(_2262_),
    .A1(net205),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6190_ (.Y(_2266_),
    .A(_2261_),
    .B(_2265_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(net165),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6192_ (.A0(rf_reg[975]),
    .A1(rf_reg[1007]),
    .S(raddr_b_i[0]),
    .X(_2268_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6193_ (.A0(rf_reg[783]),
    .A1(rf_reg[815]),
    .S(raddr_b_i[0]),
    .X(_2269_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6194_ (.Y(_2270_),
    .B1(_2269_),
    .B2(net164),
    .A2(_2268_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net165),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6196_ (.A0(rf_reg[847]),
    .A1(rf_reg[879]),
    .S(raddr_b_i[0]),
    .X(_2272_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6197_ (.A0(rf_reg[911]),
    .A1(rf_reg[943]),
    .S(raddr_b_i[0]),
    .X(_2273_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6198_ (.Y(_2274_),
    .B1(_2273_),
    .B2(net200),
    .A2(_2272_),
    .A1(net176),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6199_ (.Y(_2275_),
    .A(_2270_),
    .B(_2274_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6200_ (.Y(_2276_),
    .B1(_2275_),
    .B2(net292),
    .A2(_2266_),
    .A1(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6201_ (.B(_2258_),
    .C(_2276_),
    .A(_2249_),
    .Y(rdata_b_o[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6202_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[526]),
    .A1(rf_reg[558]),
    .A2(rf_reg[590]),
    .A3(rf_reg[622]),
    .S1(raddr_b_i[1]),
    .X(_2277_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6203_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[654]),
    .A1(rf_reg[686]),
    .A2(rf_reg[718]),
    .A3(rf_reg[750]),
    .S1(raddr_b_i[1]),
    .X(_2278_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6204_ (.Y(_2279_),
    .B1(_2278_),
    .B2(net220),
    .A2(_2277_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6205_ (.Y(_2280_),
    .A(rf_reg[46]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6206_ (.A0(rf_reg[78]),
    .A1(rf_reg[110]),
    .S(raddr_b_i[0]),
    .X(_2281_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6207_ (.Y(_2282_),
    .A(raddr_b_i[1]),
    .B(_2281_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6208_ (.B1(_2282_),
    .VDD(VDD),
    .Y(_2283_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2280_));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net165),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6210_ (.A0(rf_reg[142]),
    .A1(rf_reg[174]),
    .S(raddr_b_i[0]),
    .X(_2285_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6211_ (.A0(rf_reg[206]),
    .A1(rf_reg[238]),
    .S(raddr_b_i[0]),
    .X(_2286_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6212_ (.Y(_2287_),
    .B1(_2286_),
    .B2(net194),
    .A2(_2285_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6213_ (.A(net304),
    .B(_2287_),
    .Y(_2288_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6214_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2283_),
    .Y(_2289_),
    .B1(_2288_));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(net165),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6216_ (.A0(rf_reg[462]),
    .A1(rf_reg[494]),
    .S(raddr_b_i[0]),
    .X(_2291_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6217_ (.A0(rf_reg[334]),
    .A1(rf_reg[366]),
    .S(raddr_b_i[0]),
    .X(_2292_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6218_ (.Y(_2293_),
    .B1(_2292_),
    .B2(net175),
    .A2(_2291_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6219_ (.A0(rf_reg[398]),
    .A1(rf_reg[430]),
    .S(raddr_b_i[0]),
    .X(_2294_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6220_ (.A0(rf_reg[270]),
    .A1(rf_reg[302]),
    .S(raddr_b_i[0]),
    .X(_2295_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6221_ (.Y(_2296_),
    .B1(_2295_),
    .B2(net166),
    .A2(_2294_),
    .A1(net204),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6222_ (.Y(_2297_),
    .A(_2293_),
    .B(_2296_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6223_ (.A0(rf_reg[974]),
    .A1(rf_reg[1006]),
    .S(raddr_b_i[0]),
    .X(_2298_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(_2951_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6225_ (.A0(rf_reg[782]),
    .A1(rf_reg[814]),
    .S(raddr_b_i[0]),
    .X(_2300_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6226_ (.Y(_2301_),
    .B1(_2300_),
    .B2(net166),
    .A2(_2298_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6227_ (.A0(rf_reg[846]),
    .A1(rf_reg[878]),
    .S(raddr_b_i[0]),
    .X(_2302_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6228_ (.A0(rf_reg[910]),
    .A1(rf_reg[942]),
    .S(raddr_b_i[0]),
    .X(_2303_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6229_ (.Y(_2304_),
    .B1(_2303_),
    .B2(net204),
    .A2(_2302_),
    .A1(net175),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6230_ (.Y(_2305_),
    .A(_2301_),
    .B(_2304_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6231_ (.Y(_2306_),
    .B1(_2305_),
    .B2(net294),
    .A2(_2297_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6232_ (.B(_2289_),
    .C(_2306_),
    .A(_2279_),
    .Y(rdata_b_o[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net160),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6234_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[525]),
    .A1(rf_reg[557]),
    .A2(rf_reg[589]),
    .A3(rf_reg[621]),
    .S1(raddr_b_i[1]),
    .X(_2308_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6235_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[653]),
    .A1(rf_reg[685]),
    .A2(rf_reg[717]),
    .A3(rf_reg[749]),
    .S1(raddr_b_i[1]),
    .X(_2309_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6236_ (.Y(_2310_),
    .B1(_2309_),
    .B2(net219),
    .A2(_2308_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_2951_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout157 (.A(net158),
    .X(net157),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net158),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6240_ (.Y(_2314_),
    .A(rf_reg[45]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6241_ (.A0(rf_reg[77]),
    .A1(rf_reg[109]),
    .S(raddr_b_i[0]),
    .X(_2315_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6242_ (.Y(_2316_),
    .A(raddr_b_i[1]),
    .B(_2315_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6243_ (.B1(_2316_),
    .VDD(VDD),
    .Y(_2317_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2314_));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_3087_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6245_ (.A0(rf_reg[141]),
    .A1(rf_reg[173]),
    .S(raddr_b_i[0]),
    .X(_2319_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6246_ (.A0(rf_reg[205]),
    .A1(rf_reg[237]),
    .S(raddr_b_i[0]),
    .X(_2320_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(net155),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6248_ (.Y(_2322_),
    .B1(_2320_),
    .B2(net195),
    .A2(_2319_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6249_ (.A(net303),
    .B(_2322_),
    .Y(_2323_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6250_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2317_),
    .Y(_2324_),
    .B1(_2323_));
 sg13g2_mux2_1 _6251_ (.A0(rf_reg[461]),
    .A1(rf_reg[493]),
    .S(raddr_b_i[0]),
    .X(_2325_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6252_ (.A0(rf_reg[333]),
    .A1(rf_reg[365]),
    .S(raddr_b_i[0]),
    .X(_2326_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net154),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6254_ (.Y(_2328_),
    .B1(_2326_),
    .B2(net180),
    .A2(_2325_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6255_ (.A0(rf_reg[397]),
    .A1(rf_reg[429]),
    .S(raddr_b_i[0]),
    .X(_2329_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6256_ (.A0(rf_reg[269]),
    .A1(rf_reg[301]),
    .S(raddr_b_i[0]),
    .X(_2330_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6257_ (.Y(_2331_),
    .B1(_2330_),
    .B2(net169),
    .A2(_2329_),
    .A1(net207),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6258_ (.Y(_2332_),
    .A(_2328_),
    .B(_2331_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6259_ (.A0(rf_reg[973]),
    .A1(rf_reg[1005]),
    .S(raddr_b_i[0]),
    .X(_2333_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6260_ (.A0(rf_reg[781]),
    .A1(rf_reg[813]),
    .S(raddr_b_i[0]),
    .X(_2334_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout152 (.A(net155),
    .X(net152),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6262_ (.Y(_2336_),
    .B1(_2334_),
    .B2(net169),
    .A2(_2333_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6263_ (.A0(rf_reg[845]),
    .A1(rf_reg[877]),
    .S(raddr_b_i[0]),
    .X(_2337_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6264_ (.A0(rf_reg[909]),
    .A1(rf_reg[941]),
    .S(raddr_b_i[0]),
    .X(_2338_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6265_ (.Y(_2339_),
    .B1(_2338_),
    .B2(net207),
    .A2(_2337_),
    .A1(net180),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6266_ (.Y(_2340_),
    .A(_2336_),
    .B(_2339_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net152),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6268_ (.Y(_2342_),
    .B1(_2340_),
    .B2(net293),
    .A2(_2332_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6269_ (.B(_2324_),
    .C(_2342_),
    .A(_2310_),
    .Y(rdata_b_o[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6270_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[524]),
    .A1(rf_reg[556]),
    .A2(rf_reg[588]),
    .A3(rf_reg[620]),
    .S1(raddr_b_i[1]),
    .X(_2343_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6271_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[652]),
    .A1(rf_reg[684]),
    .A2(rf_reg[716]),
    .A3(rf_reg[748]),
    .S1(raddr_b_i[1]),
    .X(_2344_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(_3093_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6273_ (.Y(_2346_),
    .B1(_2344_),
    .B2(net218),
    .A2(_2343_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6274_ (.Y(_2347_),
    .A(rf_reg[44]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6275_ (.A0(rf_reg[76]),
    .A1(rf_reg[108]),
    .S(raddr_b_i[0]),
    .X(_2348_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6276_ (.Y(_2349_),
    .A(raddr_b_i[1]),
    .B(_2348_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6277_ (.B1(_2349_),
    .VDD(VDD),
    .Y(_2350_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2347_));
 sg13g2_mux2_1 _6278_ (.A0(rf_reg[140]),
    .A1(rf_reg[172]),
    .S(raddr_b_i[0]),
    .X(_2351_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6279_ (.A0(rf_reg[204]),
    .A1(rf_reg[236]),
    .S(raddr_b_i[0]),
    .X(_2352_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6280_ (.Y(_2353_),
    .B1(_2352_),
    .B2(net187),
    .A2(_2351_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6281_ (.A(net302),
    .B(_2353_),
    .Y(_2354_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6282_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_2350_),
    .Y(_2355_),
    .B1(_2354_));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net150),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6284_ (.A0(rf_reg[460]),
    .A1(rf_reg[492]),
    .S(raddr_b_i[0]),
    .X(_2357_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net150),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6286_ (.A0(rf_reg[332]),
    .A1(rf_reg[364]),
    .S(raddr_b_i[0]),
    .X(_2359_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6287_ (.Y(_2360_),
    .B1(_2359_),
    .B2(net175),
    .A2(_2357_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6288_ (.A0(rf_reg[396]),
    .A1(rf_reg[428]),
    .S(raddr_b_i[0]),
    .X(_2361_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6289_ (.A0(rf_reg[268]),
    .A1(rf_reg[300]),
    .S(raddr_b_i[0]),
    .X(_2362_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6290_ (.Y(_2363_),
    .B1(_2362_),
    .B2(net163),
    .A2(_2361_),
    .A1(net199),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6291_ (.Y(_2364_),
    .A(_2360_),
    .B(_2363_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6292_ (.A0(rf_reg[972]),
    .A1(rf_reg[1004]),
    .S(raddr_b_i[0]),
    .X(_2365_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6293_ (.A0(rf_reg[780]),
    .A1(rf_reg[812]),
    .S(raddr_b_i[0]),
    .X(_2366_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6294_ (.Y(_2367_),
    .B1(_2366_),
    .B2(net163),
    .A2(_2365_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6295_ (.A0(rf_reg[844]),
    .A1(rf_reg[876]),
    .S(raddr_b_i[0]),
    .X(_2368_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6296_ (.A0(rf_reg[908]),
    .A1(rf_reg[940]),
    .S(raddr_b_i[0]),
    .X(_2369_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net150),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6298_ (.Y(_2371_),
    .B1(_2369_),
    .B2(net199),
    .A2(_2368_),
    .A1(net175),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6299_ (.Y(_2372_),
    .A(_2367_),
    .B(_2371_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6300_ (.Y(_2373_),
    .B1(_2372_),
    .B2(net292),
    .A2(_2364_),
    .A1(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6301_ (.B(_2355_),
    .C(_2373_),
    .A(_2346_),
    .Y(rdata_b_o[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6302_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[541]),
    .A1(rf_reg[573]),
    .A2(rf_reg[605]),
    .A3(rf_reg[637]),
    .S1(raddr_b_i[1]),
    .X(_2374_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6303_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[669]),
    .A1(rf_reg[701]),
    .A2(rf_reg[733]),
    .A3(rf_reg[765]),
    .S1(raddr_b_i[1]),
    .X(_2375_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6304_ (.Y(_2376_),
    .B1(_2375_),
    .B2(net217),
    .A2(_2374_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6305_ (.Y(_2377_),
    .A(rf_reg[61]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6306_ (.A0(rf_reg[93]),
    .A1(rf_reg[125]),
    .S(raddr_b_i[0]),
    .X(_2378_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6307_ (.Y(_2379_),
    .A(raddr_b_i[1]),
    .B(_2378_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6308_ (.B1(_2379_),
    .VDD(VDD),
    .Y(_2380_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2377_));
 sg13g2_mux2_1 _6309_ (.A0(rf_reg[157]),
    .A1(rf_reg[189]),
    .S(raddr_b_i[0]),
    .X(_2381_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6310_ (.A0(rf_reg[221]),
    .A1(rf_reg[253]),
    .S(raddr_b_i[0]),
    .X(_2382_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6311_ (.Y(_2383_),
    .B1(_2382_),
    .B2(net186),
    .A2(_2381_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6312_ (.A(net301),
    .B(_2383_),
    .Y(_2384_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6313_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2380_),
    .Y(_2385_),
    .B1(_2384_));
 sg13g2_mux2_1 _6314_ (.A0(rf_reg[477]),
    .A1(rf_reg[509]),
    .S(raddr_b_i[0]),
    .X(_2386_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6315_ (.A0(rf_reg[349]),
    .A1(rf_reg[381]),
    .S(raddr_b_i[0]),
    .X(_2387_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6316_ (.Y(_2388_),
    .B1(_2387_),
    .B2(net172),
    .A2(_2386_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6317_ (.A0(rf_reg[413]),
    .A1(rf_reg[445]),
    .S(raddr_b_i[0]),
    .X(_2389_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6318_ (.A0(rf_reg[285]),
    .A1(rf_reg[317]),
    .S(raddr_b_i[0]),
    .X(_2390_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6319_ (.Y(_2391_),
    .B1(_2390_),
    .B2(net161),
    .A2(_2389_),
    .A1(net197),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6320_ (.Y(_2392_),
    .A(_2388_),
    .B(_2391_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6321_ (.A0(rf_reg[989]),
    .A1(rf_reg[1021]),
    .S(raddr_b_i[0]),
    .X(_2393_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6322_ (.A0(rf_reg[797]),
    .A1(rf_reg[829]),
    .S(raddr_b_i[0]),
    .X(_2394_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6323_ (.Y(_2395_),
    .B1(_2394_),
    .B2(net162),
    .A2(_2393_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6324_ (.A0(rf_reg[861]),
    .A1(rf_reg[893]),
    .S(raddr_b_i[0]),
    .X(_2396_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6325_ (.A0(rf_reg[925]),
    .A1(rf_reg[957]),
    .S(raddr_b_i[0]),
    .X(_2397_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6326_ (.Y(_2398_),
    .B1(_2397_),
    .B2(net198),
    .A2(_2396_),
    .A1(net173),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6327_ (.Y(_2399_),
    .A(_2395_),
    .B(_2398_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6328_ (.Y(_2400_),
    .B1(_2399_),
    .B2(net291),
    .A2(_2392_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6329_ (.B(_2385_),
    .C(_2400_),
    .A(_2376_),
    .Y(rdata_b_o[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6330_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[523]),
    .A1(rf_reg[555]),
    .A2(rf_reg[587]),
    .A3(rf_reg[619]),
    .S1(raddr_b_i[1]),
    .X(_2401_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6331_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[651]),
    .A1(rf_reg[683]),
    .A2(rf_reg[715]),
    .A3(rf_reg[747]),
    .S1(raddr_b_i[1]),
    .X(_2402_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6332_ (.Y(_2403_),
    .B1(_2402_),
    .B2(net220),
    .A2(_2401_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6333_ (.Y(_2404_),
    .A(rf_reg[43]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6334_ (.A0(rf_reg[75]),
    .A1(rf_reg[107]),
    .S(raddr_b_i[0]),
    .X(_2405_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6335_ (.Y(_2406_),
    .A(raddr_b_i[1]),
    .B(_2405_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6336_ (.B1(_2406_),
    .VDD(VDD),
    .Y(_2407_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2404_));
 sg13g2_mux2_1 _6337_ (.A0(rf_reg[139]),
    .A1(rf_reg[171]),
    .S(raddr_b_i[0]),
    .X(_2408_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6338_ (.A0(rf_reg[203]),
    .A1(rf_reg[235]),
    .S(raddr_b_i[0]),
    .X(_2409_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6339_ (.Y(_2410_),
    .B1(_2409_),
    .B2(net194),
    .A2(_2408_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6340_ (.A(net304),
    .B(_2410_),
    .Y(_2411_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6341_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2407_),
    .Y(_2412_),
    .B1(_2411_));
 sg13g2_mux2_1 _6342_ (.A0(rf_reg[459]),
    .A1(rf_reg[491]),
    .S(raddr_b_i[0]),
    .X(_2413_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6343_ (.A0(rf_reg[331]),
    .A1(rf_reg[363]),
    .S(raddr_b_i[0]),
    .X(_2414_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6344_ (.Y(_2415_),
    .B1(_2414_),
    .B2(net177),
    .A2(_2413_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6345_ (.A0(rf_reg[395]),
    .A1(rf_reg[427]),
    .S(raddr_b_i[0]),
    .X(_2416_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6346_ (.A0(rf_reg[267]),
    .A1(rf_reg[299]),
    .S(raddr_b_i[0]),
    .X(_2417_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6347_ (.Y(_2418_),
    .B1(_2417_),
    .B2(net166),
    .A2(_2416_),
    .A1(net204),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6348_ (.Y(_2419_),
    .A(_2415_),
    .B(_2418_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6349_ (.A0(rf_reg[971]),
    .A1(rf_reg[1003]),
    .S(raddr_b_i[0]),
    .X(_2420_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6350_ (.A0(rf_reg[779]),
    .A1(rf_reg[811]),
    .S(raddr_b_i[0]),
    .X(_2421_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6351_ (.Y(_2422_),
    .B1(_2421_),
    .B2(net166),
    .A2(_2420_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net147),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6353_ (.A0(rf_reg[843]),
    .A1(rf_reg[875]),
    .S(raddr_b_i[0]),
    .X(_2424_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(_3099_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6355_ (.A0(rf_reg[907]),
    .A1(rf_reg[939]),
    .S(raddr_b_i[0]),
    .X(_2426_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6356_ (.Y(_2427_),
    .B1(_2426_),
    .B2(net204),
    .A2(_2424_),
    .A1(net177),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6357_ (.Y(_2428_),
    .A(_2422_),
    .B(_2427_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6358_ (.Y(_2429_),
    .B1(_2428_),
    .B2(net294),
    .A2(_2419_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6359_ (.B(_2412_),
    .C(_2429_),
    .A(_2403_),
    .Y(rdata_b_o[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net145),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6361_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[522]),
    .A1(rf_reg[554]),
    .A2(rf_reg[586]),
    .A3(rf_reg[618]),
    .S1(raddr_b_i[1]),
    .X(_2431_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6362_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[650]),
    .A1(rf_reg[682]),
    .A2(rf_reg[714]),
    .A3(rf_reg[746]),
    .S1(raddr_b_i[1]),
    .X(_2432_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6363_ (.Y(_2433_),
    .B1(_2432_),
    .B2(net218),
    .A2(_2431_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6364_ (.Y(_2434_),
    .A(rf_reg[42]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6365_ (.A0(rf_reg[74]),
    .A1(rf_reg[106]),
    .S(raddr_b_i[0]),
    .X(_2435_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6366_ (.Y(_2436_),
    .A(raddr_b_i[1]),
    .B(_2435_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6367_ (.B1(_2436_),
    .VDD(VDD),
    .Y(_2437_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2434_));
 sg13g2_mux2_1 _6368_ (.A0(rf_reg[138]),
    .A1(rf_reg[170]),
    .S(raddr_b_i[0]),
    .X(_2438_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net145),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6370_ (.A0(rf_reg[202]),
    .A1(rf_reg[234]),
    .S(raddr_b_i[0]),
    .X(_2440_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6371_ (.Y(_2441_),
    .B1(_2440_),
    .B2(net187),
    .A2(_2438_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6372_ (.A(net302),
    .B(_2441_),
    .Y(_2442_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6373_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_2437_),
    .Y(_2443_),
    .B1(_2442_));
 sg13g2_mux2_1 _6374_ (.A0(rf_reg[458]),
    .A1(rf_reg[490]),
    .S(raddr_b_i[0]),
    .X(_2444_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6375_ (.A0(rf_reg[330]),
    .A1(rf_reg[362]),
    .S(raddr_b_i[0]),
    .X(_2445_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6376_ (.Y(_2446_),
    .B1(_2445_),
    .B2(net175),
    .A2(_2444_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6377_ (.A0(rf_reg[394]),
    .A1(rf_reg[426]),
    .S(raddr_b_i[0]),
    .X(_2447_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6378_ (.A0(rf_reg[266]),
    .A1(rf_reg[298]),
    .S(raddr_b_i[0]),
    .X(_2448_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6379_ (.Y(_2449_),
    .B1(_2448_),
    .B2(net163),
    .A2(_2447_),
    .A1(net199),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6380_ (.Y(_2450_),
    .A(_2446_),
    .B(_2449_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6381_ (.A0(rf_reg[970]),
    .A1(rf_reg[1002]),
    .S(raddr_b_i[0]),
    .X(_2451_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6382_ (.A0(rf_reg[778]),
    .A1(rf_reg[810]),
    .S(raddr_b_i[0]),
    .X(_2452_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6383_ (.Y(_2453_),
    .B1(_2452_),
    .B2(net164),
    .A2(_2451_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6384_ (.A0(rf_reg[842]),
    .A1(rf_reg[874]),
    .S(raddr_b_i[0]),
    .X(_2454_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6385_ (.A0(rf_reg[906]),
    .A1(rf_reg[938]),
    .S(raddr_b_i[0]),
    .X(_2455_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6386_ (.Y(_2456_),
    .B1(_2455_),
    .B2(net200),
    .A2(_2454_),
    .A1(net176),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6387_ (.Y(_2457_),
    .A(_2453_),
    .B(_2456_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6388_ (.Y(_2458_),
    .B1(_2457_),
    .B2(net292),
    .A2(_2450_),
    .A1(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6389_ (.B(_2443_),
    .C(_2458_),
    .A(_2433_),
    .Y(rdata_b_o[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6390_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[521]),
    .A1(rf_reg[553]),
    .A2(rf_reg[585]),
    .A3(rf_reg[617]),
    .S1(raddr_b_i[1]),
    .X(_2459_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6391_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[649]),
    .A1(rf_reg[681]),
    .A2(rf_reg[713]),
    .A3(rf_reg[745]),
    .S1(raddr_b_i[1]),
    .X(_2460_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6392_ (.Y(_2461_),
    .B1(_2460_),
    .B2(net217),
    .A2(_2459_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6393_ (.Y(_2462_),
    .A(rf_reg[41]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6394_ (.A0(rf_reg[73]),
    .A1(rf_reg[105]),
    .S(raddr_b_i[0]),
    .X(_2463_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6395_ (.Y(_2464_),
    .A(raddr_b_i[1]),
    .B(_2463_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6396_ (.B1(_2464_),
    .VDD(VDD),
    .Y(_2465_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2462_));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net145),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6398_ (.A0(rf_reg[137]),
    .A1(rf_reg[169]),
    .S(raddr_b_i[0]),
    .X(_2467_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6399_ (.A0(rf_reg[201]),
    .A1(rf_reg[233]),
    .S(raddr_b_i[0]),
    .X(_2468_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6400_ (.Y(_2469_),
    .B1(_2468_),
    .B2(net186),
    .A2(_2467_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6401_ (.A(net301),
    .B(_2469_),
    .Y(_2470_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6402_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2465_),
    .Y(_2471_),
    .B1(_2470_));
 sg13g2_mux2_1 _6403_ (.A0(rf_reg[457]),
    .A1(rf_reg[489]),
    .S(raddr_b_i[0]),
    .X(_2472_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6404_ (.A0(rf_reg[329]),
    .A1(rf_reg[361]),
    .S(raddr_b_i[0]),
    .X(_2473_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6405_ (.Y(_2474_),
    .B1(_2473_),
    .B2(net172),
    .A2(_2472_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net142),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6407_ (.A0(rf_reg[393]),
    .A1(rf_reg[425]),
    .S(raddr_b_i[0]),
    .X(_2476_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(_3105_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6409_ (.A0(rf_reg[265]),
    .A1(rf_reg[297]),
    .S(raddr_b_i[0]),
    .X(_2478_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6410_ (.Y(_2479_),
    .B1(_2478_),
    .B2(net161),
    .A2(_2476_),
    .A1(net197),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6411_ (.Y(_2480_),
    .A(_2474_),
    .B(_2479_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6412_ (.A0(rf_reg[969]),
    .A1(rf_reg[1001]),
    .S(raddr_b_i[0]),
    .X(_2481_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6413_ (.A0(rf_reg[777]),
    .A1(rf_reg[809]),
    .S(raddr_b_i[0]),
    .X(_2482_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6414_ (.Y(_2483_),
    .B1(_2482_),
    .B2(net161),
    .A2(_2481_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6415_ (.A0(rf_reg[841]),
    .A1(rf_reg[873]),
    .S(raddr_b_i[0]),
    .X(_2484_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6416_ (.A0(rf_reg[905]),
    .A1(rf_reg[937]),
    .S(raddr_b_i[0]),
    .X(_2485_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6417_ (.Y(_2486_),
    .B1(_2485_),
    .B2(net197),
    .A2(_2484_),
    .A1(net172),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6418_ (.Y(_2487_),
    .A(_2483_),
    .B(_2486_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6419_ (.Y(_2488_),
    .B1(_2487_),
    .B2(net291),
    .A2(_2480_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6420_ (.B(_2471_),
    .C(_2488_),
    .A(_2461_),
    .Y(rdata_b_o[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net140),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6422_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[520]),
    .A1(rf_reg[552]),
    .A2(rf_reg[584]),
    .A3(rf_reg[616]),
    .S1(raddr_b_i[1]),
    .X(_2490_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6423_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[648]),
    .A1(rf_reg[680]),
    .A2(rf_reg[712]),
    .A3(rf_reg[744]),
    .S1(raddr_b_i[1]),
    .X(_2491_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6424_ (.Y(_2492_),
    .B1(_2491_),
    .B2(net217),
    .A2(_2490_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6425_ (.Y(_2493_),
    .A(rf_reg[40]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net140),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6427_ (.A0(rf_reg[72]),
    .A1(rf_reg[104]),
    .S(raddr_b_i[0]),
    .X(_2495_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6428_ (.Y(_2496_),
    .A(raddr_b_i[1]),
    .B(_2495_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6429_ (.B1(_2496_),
    .VDD(VDD),
    .Y(_2497_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2493_));
 sg13g2_mux2_1 _6430_ (.A0(rf_reg[136]),
    .A1(rf_reg[168]),
    .S(raddr_b_i[0]),
    .X(_2498_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6431_ (.A0(rf_reg[200]),
    .A1(rf_reg[232]),
    .S(raddr_b_i[0]),
    .X(_2499_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6432_ (.Y(_2500_),
    .B1(_2499_),
    .B2(net186),
    .A2(_2498_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6433_ (.A(net302),
    .B(_2500_),
    .Y(_2501_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6434_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2497_),
    .Y(_2502_),
    .B1(_2501_));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net140),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6436_ (.A0(rf_reg[456]),
    .A1(rf_reg[488]),
    .S(raddr_b_i[0]),
    .X(_2504_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6437_ (.A0(rf_reg[328]),
    .A1(rf_reg[360]),
    .S(raddr_b_i[0]),
    .X(_2505_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6438_ (.Y(_2506_),
    .B1(_2505_),
    .B2(net172),
    .A2(_2504_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net137),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6440_ (.A0(rf_reg[392]),
    .A1(rf_reg[424]),
    .S(raddr_b_i[0]),
    .X(_2508_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6441_ (.A0(rf_reg[264]),
    .A1(rf_reg[296]),
    .S(raddr_b_i[0]),
    .X(_2509_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6442_ (.Y(_2510_),
    .B1(_2509_),
    .B2(net163),
    .A2(_2508_),
    .A1(net199),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6443_ (.Y(_2511_),
    .A(_2506_),
    .B(_2510_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6444_ (.A0(rf_reg[968]),
    .A1(rf_reg[1000]),
    .S(raddr_b_i[0]),
    .X(_2512_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6445_ (.A0(rf_reg[776]),
    .A1(rf_reg[808]),
    .S(raddr_b_i[0]),
    .X(_2513_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6446_ (.Y(_2514_),
    .B1(_2513_),
    .B2(net163),
    .A2(_2512_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6447_ (.A0(rf_reg[840]),
    .A1(rf_reg[872]),
    .S(raddr_b_i[0]),
    .X(_2515_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6448_ (.A0(rf_reg[904]),
    .A1(rf_reg[936]),
    .S(raddr_b_i[0]),
    .X(_2516_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6449_ (.Y(_2517_),
    .B1(_2516_),
    .B2(net199),
    .A2(_2515_),
    .A1(net172),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6450_ (.Y(_2518_),
    .A(_2514_),
    .B(_2517_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6451_ (.Y(_2519_),
    .B1(_2518_),
    .B2(net291),
    .A2(_2511_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6452_ (.B(_2502_),
    .C(_2519_),
    .A(_2492_),
    .Y(rdata_b_o[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6453_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[519]),
    .A1(rf_reg[551]),
    .A2(rf_reg[583]),
    .A3(rf_reg[615]),
    .S1(raddr_b_i[1]),
    .X(_2520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6454_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[647]),
    .A1(rf_reg[679]),
    .A2(rf_reg[711]),
    .A3(rf_reg[743]),
    .S1(raddr_b_i[1]),
    .X(_2521_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6455_ (.Y(_2522_),
    .B1(_2521_),
    .B2(net219),
    .A2(_2520_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6456_ (.Y(_2523_),
    .A(rf_reg[39]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_3133_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6458_ (.A0(rf_reg[71]),
    .A1(rf_reg[103]),
    .S(raddr_b_i[0]),
    .X(_2525_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6459_ (.Y(_2526_),
    .A(raddr_b_i[1]),
    .B(_2525_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6460_ (.B1(_2526_),
    .VDD(VDD),
    .Y(_2527_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2523_));
 sg13g2_mux2_1 _6461_ (.A0(rf_reg[135]),
    .A1(rf_reg[167]),
    .S(raddr_b_i[0]),
    .X(_2528_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6462_ (.A0(rf_reg[199]),
    .A1(rf_reg[231]),
    .S(raddr_b_i[0]),
    .X(_2529_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6463_ (.Y(_2530_),
    .B1(_2529_),
    .B2(net195),
    .A2(_2528_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6464_ (.A(net303),
    .B(_2530_),
    .Y(_2531_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6465_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2527_),
    .Y(_2532_),
    .B1(_2531_));
 sg13g2_mux2_1 _6466_ (.A0(rf_reg[455]),
    .A1(rf_reg[487]),
    .S(raddr_b_i[0]),
    .X(_2533_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6467_ (.A0(rf_reg[327]),
    .A1(rf_reg[359]),
    .S(raddr_b_i[0]),
    .X(_2534_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6468_ (.Y(_2535_),
    .B1(_2534_),
    .B2(net179),
    .A2(_2533_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6469_ (.A0(rf_reg[391]),
    .A1(rf_reg[423]),
    .S(raddr_b_i[0]),
    .X(_2536_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6470_ (.A0(rf_reg[263]),
    .A1(rf_reg[295]),
    .S(raddr_b_i[0]),
    .X(_2537_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6471_ (.Y(_2538_),
    .B1(_2537_),
    .B2(net168),
    .A2(_2536_),
    .A1(net206),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6472_ (.Y(_2539_),
    .A(_2535_),
    .B(_2538_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net135),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6474_ (.A0(rf_reg[967]),
    .A1(rf_reg[999]),
    .S(raddr_b_i[0]),
    .X(_2541_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6475_ (.A0(rf_reg[775]),
    .A1(rf_reg[807]),
    .S(raddr_b_i[0]),
    .X(_2542_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6476_ (.Y(_2543_),
    .B1(_2542_),
    .B2(net168),
    .A2(_2541_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6477_ (.A0(rf_reg[839]),
    .A1(rf_reg[871]),
    .S(raddr_b_i[0]),
    .X(_2544_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6478_ (.A0(rf_reg[903]),
    .A1(rf_reg[935]),
    .S(raddr_b_i[0]),
    .X(_2545_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6479_ (.Y(_2546_),
    .B1(_2545_),
    .B2(net206),
    .A2(_2544_),
    .A1(net179),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6480_ (.Y(_2547_),
    .A(_2543_),
    .B(_2546_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6481_ (.Y(_2548_),
    .B1(_2547_),
    .B2(net293),
    .A2(_2539_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6482_ (.B(_2532_),
    .C(_2548_),
    .A(_2522_),
    .Y(rdata_b_o[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6483_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[518]),
    .A1(rf_reg[550]),
    .A2(rf_reg[582]),
    .A3(rf_reg[614]),
    .S1(raddr_b_i[1]),
    .X(_2549_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net135),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net135),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6486_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[646]),
    .A1(rf_reg[678]),
    .A2(rf_reg[710]),
    .A3(rf_reg[742]),
    .S1(raddr_b_i[1]),
    .X(_2552_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6487_ (.Y(_2553_),
    .B1(_2552_),
    .B2(net218),
    .A2(_2549_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6488_ (.Y(_2554_),
    .A(rf_reg[38]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6489_ (.A0(rf_reg[70]),
    .A1(rf_reg[102]),
    .S(raddr_b_i[0]),
    .X(_2555_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6490_ (.Y(_2556_),
    .A(raddr_b_i[1]),
    .B(_2555_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6491_ (.B1(_2556_),
    .VDD(VDD),
    .Y(_2557_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2554_));
 sg13g2_mux2_1 _6492_ (.A0(rf_reg[134]),
    .A1(rf_reg[166]),
    .S(raddr_b_i[0]),
    .X(_2558_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6493_ (.A0(rf_reg[198]),
    .A1(rf_reg[230]),
    .S(raddr_b_i[0]),
    .X(_2559_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6494_ (.Y(_2560_),
    .B1(_2559_),
    .B2(net187),
    .A2(_2558_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6495_ (.A(net301),
    .B(_2560_),
    .Y(_2561_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6496_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2557_),
    .Y(_2562_),
    .B1(_2561_));
 sg13g2_mux2_1 _6497_ (.A0(rf_reg[454]),
    .A1(rf_reg[486]),
    .S(raddr_b_i[0]),
    .X(_2563_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6498_ (.A0(rf_reg[326]),
    .A1(rf_reg[358]),
    .S(raddr_b_i[0]),
    .X(_2564_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6499_ (.Y(_2565_),
    .B1(_2564_),
    .B2(net176),
    .A2(_2563_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6500_ (.A0(rf_reg[390]),
    .A1(rf_reg[422]),
    .S(raddr_b_i[0]),
    .X(_2566_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6501_ (.A0(rf_reg[262]),
    .A1(rf_reg[294]),
    .S(raddr_b_i[0]),
    .X(_2567_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net132),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6503_ (.Y(_2569_),
    .B1(_2567_),
    .B2(net164),
    .A2(_2566_),
    .A1(net200),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6504_ (.Y(_2570_),
    .A(_2565_),
    .B(_2569_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_3143_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6506_ (.A0(rf_reg[966]),
    .A1(rf_reg[998]),
    .S(raddr_b_i[0]),
    .X(_2572_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6507_ (.A0(rf_reg[774]),
    .A1(rf_reg[806]),
    .S(raddr_b_i[0]),
    .X(_2573_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6508_ (.Y(_2574_),
    .B1(_2573_),
    .B2(net164),
    .A2(_2572_),
    .A1(net185),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net130),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6510_ (.A0(rf_reg[838]),
    .A1(rf_reg[870]),
    .S(raddr_b_i[0]),
    .X(_2576_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6511_ (.A0(rf_reg[902]),
    .A1(rf_reg[934]),
    .S(raddr_b_i[0]),
    .X(_2577_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6512_ (.Y(_2578_),
    .B1(_2577_),
    .B2(net200),
    .A2(_2576_),
    .A1(net174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6513_ (.Y(_2579_),
    .A(_2574_),
    .B(_2578_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6514_ (.Y(_2580_),
    .B1(_2579_),
    .B2(net292),
    .A2(_2570_),
    .A1(net297),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6515_ (.B(_2562_),
    .C(_2580_),
    .A(_2553_),
    .Y(rdata_b_o[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6516_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[517]),
    .A1(rf_reg[549]),
    .A2(rf_reg[581]),
    .A3(rf_reg[613]),
    .S1(raddr_b_i[1]),
    .X(_2581_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6517_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[645]),
    .A1(rf_reg[677]),
    .A2(rf_reg[709]),
    .A3(rf_reg[741]),
    .S1(raddr_b_i[1]),
    .X(_2582_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6518_ (.Y(_2583_),
    .B1(_2582_),
    .B2(net219),
    .A2(_2581_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6519_ (.Y(_2584_),
    .A(rf_reg[37]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6520_ (.A0(rf_reg[69]),
    .A1(rf_reg[101]),
    .S(raddr_b_i[0]),
    .X(_2585_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6521_ (.Y(_2586_),
    .A(raddr_b_i[1]),
    .B(_2585_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6522_ (.B1(_2586_),
    .VDD(VDD),
    .Y(_2587_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2584_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net129),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6524_ (.A0(rf_reg[133]),
    .A1(rf_reg[165]),
    .S(raddr_b_i[0]),
    .X(_2589_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6525_ (.A0(rf_reg[197]),
    .A1(rf_reg[229]),
    .S(raddr_b_i[0]),
    .X(_2590_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6526_ (.Y(_2591_),
    .B1(_2590_),
    .B2(net195),
    .A2(_2589_),
    .A1(net211),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6527_ (.A(net303),
    .B(_2591_),
    .Y(_2592_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6528_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2587_),
    .Y(_2593_),
    .B1(_2592_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net130),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6530_ (.A0(rf_reg[453]),
    .A1(rf_reg[485]),
    .S(raddr_b_i[0]),
    .X(_2595_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6531_ (.A0(rf_reg[325]),
    .A1(rf_reg[357]),
    .S(raddr_b_i[0]),
    .X(_2596_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6532_ (.Y(_2597_),
    .B1(_2596_),
    .B2(net179),
    .A2(_2595_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6533_ (.A0(rf_reg[389]),
    .A1(rf_reg[421]),
    .S(raddr_b_i[0]),
    .X(_2598_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6534_ (.A0(rf_reg[261]),
    .A1(rf_reg[293]),
    .S(raddr_b_i[0]),
    .X(_2599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6535_ (.Y(_2600_),
    .B1(_2599_),
    .B2(net170),
    .A2(_2598_),
    .A1(net206),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6536_ (.Y(_2601_),
    .A(_2597_),
    .B(_2600_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6537_ (.A0(rf_reg[965]),
    .A1(rf_reg[997]),
    .S(raddr_b_i[0]),
    .X(_2602_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(net130),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6539_ (.A0(rf_reg[773]),
    .A1(rf_reg[805]),
    .S(raddr_b_i[0]),
    .X(_2604_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6540_ (.Y(_2605_),
    .B1(_2604_),
    .B2(net168),
    .A2(_2602_),
    .A1(net193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6541_ (.A0(rf_reg[837]),
    .A1(rf_reg[869]),
    .S(raddr_b_i[0]),
    .X(_2606_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6542_ (.A0(rf_reg[901]),
    .A1(rf_reg[933]),
    .S(raddr_b_i[0]),
    .X(_2607_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6543_ (.Y(_2608_),
    .B1(_2607_),
    .B2(net206),
    .A2(_2606_),
    .A1(net179),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6544_ (.Y(_2609_),
    .A(_2605_),
    .B(_2608_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6545_ (.Y(_2610_),
    .B1(_2609_),
    .B2(net293),
    .A2(_2601_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6546_ (.B(_2593_),
    .C(_2610_),
    .A(_2583_),
    .Y(rdata_b_o[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_3148_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6548_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[516]),
    .A1(rf_reg[548]),
    .A2(rf_reg[580]),
    .A3(rf_reg[612]),
    .S1(raddr_b_i[1]),
    .X(_2612_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6549_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[644]),
    .A1(rf_reg[676]),
    .A2(rf_reg[708]),
    .A3(rf_reg[740]),
    .S1(raddr_b_i[1]),
    .X(_2613_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6550_ (.Y(_2614_),
    .B1(_2613_),
    .B2(net217),
    .A2(_2612_),
    .A1(net223),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net125),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(net124),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net125),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6554_ (.Y(_2618_),
    .A(rf_reg[36]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6555_ (.A0(rf_reg[68]),
    .A1(rf_reg[100]),
    .S(raddr_b_i[0]),
    .X(_2619_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6556_ (.Y(_2620_),
    .A(raddr_b_i[1]),
    .B(_2619_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6557_ (.B1(_2620_),
    .VDD(VDD),
    .Y(_2621_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2618_));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net122),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6559_ (.A0(rf_reg[132]),
    .A1(rf_reg[164]),
    .S(raddr_b_i[0]),
    .X(_2623_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6560_ (.A0(rf_reg[196]),
    .A1(rf_reg[228]),
    .S(raddr_b_i[0]),
    .X(_2624_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_3153_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6562_ (.Y(_2626_),
    .B1(_2624_),
    .B2(net186),
    .A2(_2623_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6563_ (.A(net301),
    .B(_2626_),
    .Y(_2627_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6564_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_2621_),
    .Y(_2628_),
    .B1(_2627_));
 sg13g2_mux2_1 _6565_ (.A0(rf_reg[452]),
    .A1(rf_reg[484]),
    .S(raddr_b_i[0]),
    .X(_2629_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6566_ (.A0(rf_reg[324]),
    .A1(rf_reg[356]),
    .S(raddr_b_i[0]),
    .X(_2630_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(net120),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6568_ (.Y(_2632_),
    .B1(_2630_),
    .B2(net172),
    .A2(_2629_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6569_ (.A0(rf_reg[388]),
    .A1(rf_reg[420]),
    .S(raddr_b_i[0]),
    .X(_2633_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6570_ (.A0(rf_reg[260]),
    .A1(rf_reg[292]),
    .S(raddr_b_i[0]),
    .X(_2634_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6571_ (.Y(_2635_),
    .B1(_2634_),
    .B2(net161),
    .A2(_2633_),
    .A1(net197),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6572_ (.Y(_2636_),
    .A(_2632_),
    .B(_2635_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6573_ (.A0(rf_reg[964]),
    .A1(rf_reg[996]),
    .S(raddr_b_i[0]),
    .X(_2637_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6574_ (.A0(rf_reg[772]),
    .A1(rf_reg[804]),
    .S(raddr_b_i[0]),
    .X(_2638_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(net119),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6576_ (.Y(_2640_),
    .B1(_2638_),
    .B2(net162),
    .A2(_2637_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6577_ (.A0(rf_reg[836]),
    .A1(rf_reg[868]),
    .S(raddr_b_i[0]),
    .X(_2641_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6578_ (.A0(rf_reg[900]),
    .A1(rf_reg[932]),
    .S(raddr_b_i[0]),
    .X(_2642_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6579_ (.Y(_2643_),
    .B1(_2642_),
    .B2(net198),
    .A2(_2641_),
    .A1(net173),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6580_ (.Y(_2644_),
    .A(_2640_),
    .B(_2643_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(net120),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6582_ (.Y(_2646_),
    .B1(_2644_),
    .B2(net291),
    .A2(_2636_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6583_ (.B(_2628_),
    .C(_2646_),
    .A(_2614_),
    .Y(rdata_b_o[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6584_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[515]),
    .A1(rf_reg[547]),
    .A2(rf_reg[579]),
    .A3(rf_reg[611]),
    .S1(raddr_b_i[1]),
    .X(_2647_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6585_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[643]),
    .A1(rf_reg[675]),
    .A2(rf_reg[707]),
    .A3(rf_reg[739]),
    .S1(raddr_b_i[1]),
    .X(_2648_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(net120),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6587_ (.Y(_2650_),
    .B1(_2648_),
    .B2(net220),
    .A2(_2647_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6588_ (.Y(_2651_),
    .A(rf_reg[35]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6589_ (.A0(rf_reg[67]),
    .A1(rf_reg[99]),
    .S(raddr_b_i[0]),
    .X(_2652_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6590_ (.Y(_2653_),
    .A(raddr_b_i[1]),
    .B(_2652_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6591_ (.B1(_2653_),
    .VDD(VDD),
    .Y(_2654_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2651_));
 sg13g2_mux2_1 _6592_ (.A0(rf_reg[131]),
    .A1(rf_reg[163]),
    .S(raddr_b_i[0]),
    .X(_2655_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6593_ (.A0(rf_reg[195]),
    .A1(rf_reg[227]),
    .S(raddr_b_i[0]),
    .X(_2656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6594_ (.Y(_2657_),
    .B1(_2656_),
    .B2(net195),
    .A2(_2655_),
    .A1(net211),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6595_ (.A(net305),
    .B(_2657_),
    .Y(_2658_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6596_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2654_),
    .Y(_2659_),
    .B1(_2658_));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_3157_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6598_ (.A0(rf_reg[451]),
    .A1(rf_reg[483]),
    .S(raddr_b_i[0]),
    .X(_2661_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6600_ (.A0(rf_reg[323]),
    .A1(rf_reg[355]),
    .S(raddr_b_i[0]),
    .X(_2663_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6601_ (.Y(_2664_),
    .B1(_2663_),
    .B2(net181),
    .A2(_2661_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6602_ (.A0(rf_reg[387]),
    .A1(rf_reg[419]),
    .S(raddr_b_i[0]),
    .X(_2665_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6603_ (.A0(rf_reg[259]),
    .A1(rf_reg[291]),
    .S(raddr_b_i[0]),
    .X(_2666_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6604_ (.Y(_2667_),
    .B1(_2666_),
    .B2(net170),
    .A2(_2665_),
    .A1(net206),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6605_ (.Y(_2668_),
    .A(_2664_),
    .B(_2667_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6606_ (.A0(rf_reg[963]),
    .A1(rf_reg[995]),
    .S(raddr_b_i[0]),
    .X(_2669_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6607_ (.A0(rf_reg[771]),
    .A1(rf_reg[803]),
    .S(raddr_b_i[0]),
    .X(_2670_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6608_ (.Y(_2671_),
    .B1(_2670_),
    .B2(net170),
    .A2(_2669_),
    .A1(net193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6609_ (.A0(rf_reg[835]),
    .A1(rf_reg[867]),
    .S(raddr_b_i[0]),
    .X(_2672_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6610_ (.A0(rf_reg[899]),
    .A1(rf_reg[931]),
    .S(raddr_b_i[0]),
    .X(_2673_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(net114),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6612_ (.Y(_2675_),
    .B1(_2673_),
    .B2(net208),
    .A2(_2672_),
    .A1(net179),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6613_ (.Y(_2676_),
    .A(_2671_),
    .B(_2675_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6614_ (.Y(_2677_),
    .B1(_2676_),
    .B2(net294),
    .A2(_2668_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6615_ (.B(_2659_),
    .C(_2677_),
    .A(_2650_),
    .Y(rdata_b_o[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6616_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[514]),
    .A1(rf_reg[546]),
    .A2(rf_reg[578]),
    .A3(rf_reg[610]),
    .S1(raddr_b_i[1]),
    .X(_2678_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6617_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[642]),
    .A1(rf_reg[674]),
    .A2(rf_reg[706]),
    .A3(rf_reg[738]),
    .S1(raddr_b_i[1]),
    .X(_2679_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6618_ (.Y(_2680_),
    .B1(_2679_),
    .B2(net217),
    .A2(_2678_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6619_ (.Y(_2681_),
    .A(rf_reg[34]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6620_ (.A0(rf_reg[66]),
    .A1(rf_reg[98]),
    .S(raddr_b_i[0]),
    .X(_2682_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6621_ (.Y(_2683_),
    .A(raddr_b_i[1]),
    .B(_2682_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6622_ (.B1(_2683_),
    .VDD(VDD),
    .Y(_2684_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2681_));
 sg13g2_mux2_1 _6623_ (.A0(rf_reg[130]),
    .A1(rf_reg[162]),
    .S(raddr_b_i[0]),
    .X(_2685_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6624_ (.A0(rf_reg[194]),
    .A1(rf_reg[226]),
    .S(raddr_b_i[0]),
    .X(_2686_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6625_ (.Y(_2687_),
    .B1(_2686_),
    .B2(net187),
    .A2(_2685_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6626_ (.A(net301),
    .B(_2687_),
    .Y(_2688_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6627_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2684_),
    .Y(_2689_),
    .B1(_2688_));
 sg13g2_mux2_1 _6628_ (.A0(rf_reg[450]),
    .A1(rf_reg[482]),
    .S(raddr_b_i[0]),
    .X(_2690_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6629_ (.A0(rf_reg[322]),
    .A1(rf_reg[354]),
    .S(raddr_b_i[0]),
    .X(_2691_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6630_ (.Y(_2692_),
    .B1(_2691_),
    .B2(net172),
    .A2(_2690_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6631_ (.A0(rf_reg[386]),
    .A1(rf_reg[418]),
    .S(raddr_b_i[0]),
    .X(_2693_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6632_ (.A0(rf_reg[258]),
    .A1(rf_reg[290]),
    .S(raddr_b_i[0]),
    .X(_2694_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6633_ (.Y(_2695_),
    .B1(_2694_),
    .B2(net161),
    .A2(_2693_),
    .A1(net197),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6634_ (.Y(_2696_),
    .A(_2692_),
    .B(_2695_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6635_ (.A0(rf_reg[962]),
    .A1(rf_reg[994]),
    .S(raddr_b_i[0]),
    .X(_2697_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6636_ (.A0(rf_reg[770]),
    .A1(rf_reg[802]),
    .S(raddr_b_i[0]),
    .X(_2698_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6637_ (.Y(_2699_),
    .B1(_2698_),
    .B2(net161),
    .A2(_2697_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6638_ (.A0(rf_reg[834]),
    .A1(rf_reg[866]),
    .S(raddr_b_i[0]),
    .X(_2700_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6639_ (.A0(rf_reg[898]),
    .A1(rf_reg[930]),
    .S(raddr_b_i[0]),
    .X(_2701_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6640_ (.Y(_2702_),
    .B1(_2701_),
    .B2(net197),
    .A2(_2700_),
    .A1(net172),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6641_ (.Y(_2703_),
    .A(_2699_),
    .B(_2702_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6642_ (.Y(_2704_),
    .B1(_2703_),
    .B2(net291),
    .A2(_2696_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6643_ (.B(_2689_),
    .C(_2704_),
    .A(_2680_),
    .Y(rdata_b_o[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6644_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[540]),
    .A1(rf_reg[572]),
    .A2(rf_reg[604]),
    .A3(rf_reg[636]),
    .S1(raddr_b_i[1]),
    .X(_2705_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6645_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[668]),
    .A1(rf_reg[700]),
    .A2(rf_reg[732]),
    .A3(rf_reg[764]),
    .S1(raddr_b_i[1]),
    .X(_2706_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6646_ (.Y(_2707_),
    .B1(_2706_),
    .B2(net221),
    .A2(_2705_),
    .A1(net226),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6647_ (.Y(_2708_),
    .A(rf_reg[60]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6648_ (.A0(rf_reg[92]),
    .A1(rf_reg[124]),
    .S(raddr_b_i[0]),
    .X(_2709_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6649_ (.Y(_2710_),
    .A(raddr_b_i[1]),
    .B(_2709_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6650_ (.B1(_2710_),
    .VDD(VDD),
    .Y(_2711_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2708_));
 sg13g2_mux2_1 _6651_ (.A0(rf_reg[156]),
    .A1(rf_reg[188]),
    .S(raddr_b_i[0]),
    .X(_2712_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6652_ (.A0(rf_reg[220]),
    .A1(rf_reg[252]),
    .S(raddr_b_i[0]),
    .X(_2713_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6653_ (.Y(_2714_),
    .B1(_2713_),
    .B2(net195),
    .A2(_2712_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6654_ (.A(net305),
    .B(_2714_),
    .Y(_2715_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6655_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net216),
    .A2(_2711_),
    .Y(_2716_),
    .B1(_2715_));
 sg13g2_mux2_1 _6656_ (.A0(rf_reg[476]),
    .A1(rf_reg[508]),
    .S(raddr_b_i[0]),
    .X(_2717_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6657_ (.A0(rf_reg[348]),
    .A1(rf_reg[380]),
    .S(raddr_b_i[0]),
    .X(_2718_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6658_ (.Y(_2719_),
    .B1(_2718_),
    .B2(net180),
    .A2(_2717_),
    .A1(net193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6659_ (.A0(rf_reg[412]),
    .A1(rf_reg[444]),
    .S(raddr_b_i[0]),
    .X(_2720_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6660_ (.A0(rf_reg[284]),
    .A1(rf_reg[316]),
    .S(raddr_b_i[0]),
    .X(_2721_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6661_ (.Y(_2722_),
    .B1(_2721_),
    .B2(net169),
    .A2(_2720_),
    .A1(net207),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6662_ (.Y(_2723_),
    .A(_2719_),
    .B(_2722_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6663_ (.A0(rf_reg[988]),
    .A1(rf_reg[1020]),
    .S(raddr_b_i[0]),
    .X(_2724_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6664_ (.A0(rf_reg[796]),
    .A1(rf_reg[828]),
    .S(raddr_b_i[0]),
    .X(_2725_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6665_ (.Y(_2726_),
    .B1(_2725_),
    .B2(net169),
    .A2(_2724_),
    .A1(net193),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6666_ (.A0(rf_reg[860]),
    .A1(rf_reg[892]),
    .S(raddr_b_i[0]),
    .X(_2727_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6667_ (.A0(rf_reg[924]),
    .A1(rf_reg[956]),
    .S(raddr_b_i[0]),
    .X(_2728_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6668_ (.Y(_2729_),
    .B1(_2728_),
    .B2(net207),
    .A2(_2727_),
    .A1(net180),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6669_ (.Y(_2730_),
    .A(_2726_),
    .B(_2729_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6670_ (.Y(_2731_),
    .B1(_2730_),
    .B2(net293),
    .A2(_2723_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6671_ (.B(_2716_),
    .C(_2731_),
    .A(_2707_),
    .Y(rdata_b_o[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6672_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[513]),
    .A1(rf_reg[545]),
    .A2(rf_reg[577]),
    .A3(rf_reg[609]),
    .S1(raddr_b_i[1]),
    .X(_2732_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6673_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[641]),
    .A1(rf_reg[673]),
    .A2(rf_reg[705]),
    .A3(rf_reg[737]),
    .S1(raddr_b_i[1]),
    .X(_2733_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6674_ (.Y(_2734_),
    .B1(_2733_),
    .B2(net220),
    .A2(_2732_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6675_ (.Y(_2735_),
    .A(rf_reg[33]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6676_ (.A0(rf_reg[65]),
    .A1(rf_reg[97]),
    .S(raddr_b_i[0]),
    .X(_2736_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6677_ (.Y(_2737_),
    .A(raddr_b_i[1]),
    .B(_2736_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6678_ (.B1(_2737_),
    .VDD(VDD),
    .Y(_2738_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2735_));
 sg13g2_mux2_1 _6679_ (.A0(rf_reg[129]),
    .A1(rf_reg[161]),
    .S(raddr_b_i[0]),
    .X(_2739_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6680_ (.A0(rf_reg[193]),
    .A1(rf_reg[225]),
    .S(raddr_b_i[0]),
    .X(_2740_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6681_ (.Y(_2741_),
    .B1(_2740_),
    .B2(net194),
    .A2(_2739_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6682_ (.A(net304),
    .B(_2741_),
    .Y(_2742_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6683_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2738_),
    .Y(_2743_),
    .B1(_2742_));
 sg13g2_mux2_1 _6684_ (.A0(rf_reg[449]),
    .A1(rf_reg[481]),
    .S(raddr_b_i[0]),
    .X(_2744_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6685_ (.A0(rf_reg[321]),
    .A1(rf_reg[353]),
    .S(raddr_b_i[0]),
    .X(_2745_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6686_ (.Y(_2746_),
    .B1(_2745_),
    .B2(net177),
    .A2(_2744_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6687_ (.A0(rf_reg[385]),
    .A1(rf_reg[417]),
    .S(raddr_b_i[0]),
    .X(_2747_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6688_ (.A0(rf_reg[257]),
    .A1(rf_reg[289]),
    .S(raddr_b_i[0]),
    .X(_2748_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6689_ (.Y(_2749_),
    .B1(_2748_),
    .B2(net166),
    .A2(_2747_),
    .A1(net205),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6690_ (.Y(_2750_),
    .A(_2746_),
    .B(_2749_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6691_ (.A0(rf_reg[961]),
    .A1(rf_reg[993]),
    .S(raddr_b_i[0]),
    .X(_2751_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6692_ (.A0(rf_reg[769]),
    .A1(rf_reg[801]),
    .S(raddr_b_i[0]),
    .X(_2752_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6693_ (.Y(_2753_),
    .B1(_2752_),
    .B2(net167),
    .A2(_2751_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6694_ (.A0(rf_reg[833]),
    .A1(rf_reg[865]),
    .S(raddr_b_i[0]),
    .X(_2754_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6695_ (.A0(rf_reg[897]),
    .A1(rf_reg[929]),
    .S(raddr_b_i[0]),
    .X(_2755_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6696_ (.Y(_2756_),
    .B1(_2755_),
    .B2(net204),
    .A2(_2754_),
    .A1(net177),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6697_ (.Y(_2757_),
    .A(_2753_),
    .B(_2756_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6698_ (.Y(_2758_),
    .B1(_2757_),
    .B2(net294),
    .A2(_2750_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6699_ (.B(_2743_),
    .C(_2758_),
    .A(_2734_),
    .Y(rdata_b_o[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6700_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[512]),
    .A1(rf_reg[544]),
    .A2(rf_reg[576]),
    .A3(rf_reg[608]),
    .S1(raddr_b_i[1]),
    .X(_2759_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6701_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[640]),
    .A1(rf_reg[672]),
    .A2(rf_reg[704]),
    .A3(rf_reg[736]),
    .S1(raddr_b_i[1]),
    .X(_2760_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6702_ (.Y(_2761_),
    .B1(_2760_),
    .B2(net220),
    .A2(_2759_),
    .A1(net225),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6703_ (.Y(_2762_),
    .A(rf_reg[32]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6704_ (.A0(rf_reg[64]),
    .A1(rf_reg[96]),
    .S(raddr_b_i[0]),
    .X(_2763_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6705_ (.Y(_2764_),
    .A(raddr_b_i[1]),
    .B(_2763_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6706_ (.B1(_2764_),
    .VDD(VDD),
    .Y(_2765_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2762_));
 sg13g2_mux2_1 _6707_ (.A0(rf_reg[128]),
    .A1(rf_reg[160]),
    .S(raddr_b_i[0]),
    .X(_2766_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6708_ (.A0(rf_reg[192]),
    .A1(rf_reg[224]),
    .S(raddr_b_i[0]),
    .X(_2767_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6709_ (.Y(_2768_),
    .B1(_2767_),
    .B2(net194),
    .A2(_2766_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6710_ (.A(net304),
    .B(_2768_),
    .Y(_2769_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6711_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net215),
    .A2(_2765_),
    .Y(_2770_),
    .B1(_2769_));
 sg13g2_mux2_1 _6712_ (.A0(rf_reg[448]),
    .A1(rf_reg[480]),
    .S(raddr_b_i[0]),
    .X(_2771_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6713_ (.A0(rf_reg[320]),
    .A1(rf_reg[352]),
    .S(raddr_b_i[0]),
    .X(_2772_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6714_ (.Y(_2773_),
    .B1(_2772_),
    .B2(net177),
    .A2(_2771_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6715_ (.A0(rf_reg[384]),
    .A1(rf_reg[416]),
    .S(raddr_b_i[0]),
    .X(_2774_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6716_ (.A0(rf_reg[256]),
    .A1(rf_reg[288]),
    .S(raddr_b_i[0]),
    .X(_2775_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6717_ (.Y(_2776_),
    .B1(_2775_),
    .B2(net166),
    .A2(_2774_),
    .A1(net204),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6718_ (.Y(_2777_),
    .A(_2773_),
    .B(_2776_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6719_ (.A0(rf_reg[960]),
    .A1(rf_reg[992]),
    .S(raddr_b_i[0]),
    .X(_2778_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6720_ (.A0(rf_reg[768]),
    .A1(rf_reg[800]),
    .S(raddr_b_i[0]),
    .X(_2779_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6721_ (.Y(_2780_),
    .B1(_2779_),
    .B2(net166),
    .A2(_2778_),
    .A1(net189),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6722_ (.A0(rf_reg[832]),
    .A1(rf_reg[864]),
    .S(raddr_b_i[0]),
    .X(_2781_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6723_ (.A0(rf_reg[896]),
    .A1(rf_reg[928]),
    .S(raddr_b_i[0]),
    .X(_2782_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6724_ (.Y(_2783_),
    .B1(_2782_),
    .B2(net205),
    .A2(_2781_),
    .A1(net177),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6725_ (.Y(_2784_),
    .A(_2780_),
    .B(_2783_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6726_ (.Y(_2785_),
    .B1(_2784_),
    .B2(net294),
    .A2(_2777_),
    .A1(net299),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6727_ (.B(_2770_),
    .C(_2785_),
    .A(_2761_),
    .Y(rdata_b_o[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6728_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[539]),
    .A1(rf_reg[571]),
    .A2(rf_reg[603]),
    .A3(rf_reg[635]),
    .S1(raddr_b_i[1]),
    .X(_2786_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6729_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[667]),
    .A1(rf_reg[699]),
    .A2(rf_reg[731]),
    .A3(rf_reg[763]),
    .S1(raddr_b_i[1]),
    .X(_2787_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6730_ (.Y(_2788_),
    .B1(_2787_),
    .B2(net219),
    .A2(_2786_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6731_ (.Y(_2789_),
    .A(rf_reg[59]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6732_ (.A0(rf_reg[91]),
    .A1(rf_reg[123]),
    .S(raddr_b_i[0]),
    .X(_2790_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6733_ (.Y(_2791_),
    .A(raddr_b_i[1]),
    .B(_2790_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6734_ (.B1(_2791_),
    .VDD(VDD),
    .Y(_2792_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2789_));
 sg13g2_mux2_1 _6735_ (.A0(rf_reg[155]),
    .A1(rf_reg[187]),
    .S(raddr_b_i[0]),
    .X(_2793_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6736_ (.A0(rf_reg[219]),
    .A1(rf_reg[251]),
    .S(raddr_b_i[0]),
    .X(_2794_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6737_ (.Y(_2795_),
    .B1(_2794_),
    .B2(net194),
    .A2(_2793_),
    .A1(net209),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6738_ (.A(net303),
    .B(_2795_),
    .Y(_2796_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6739_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2792_),
    .Y(_2797_),
    .B1(_2796_));
 sg13g2_mux2_1 _6740_ (.A0(rf_reg[475]),
    .A1(rf_reg[507]),
    .S(raddr_b_i[0]),
    .X(_2798_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6741_ (.A0(rf_reg[347]),
    .A1(rf_reg[379]),
    .S(raddr_b_i[0]),
    .X(_2799_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6742_ (.Y(_2800_),
    .B1(_2799_),
    .B2(net179),
    .A2(_2798_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6743_ (.A0(rf_reg[411]),
    .A1(rf_reg[443]),
    .S(raddr_b_i[0]),
    .X(_2801_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6744_ (.A0(rf_reg[283]),
    .A1(rf_reg[315]),
    .S(raddr_b_i[0]),
    .X(_2802_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6745_ (.Y(_2803_),
    .B1(_2802_),
    .B2(net168),
    .A2(_2801_),
    .A1(net206),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6746_ (.Y(_2804_),
    .A(_2800_),
    .B(_2803_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6747_ (.A0(rf_reg[987]),
    .A1(rf_reg[1019]),
    .S(raddr_b_i[0]),
    .X(_2805_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6748_ (.A0(rf_reg[795]),
    .A1(rf_reg[827]),
    .S(raddr_b_i[0]),
    .X(_2806_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6749_ (.Y(_2807_),
    .B1(_2806_),
    .B2(net168),
    .A2(_2805_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6750_ (.A0(rf_reg[859]),
    .A1(rf_reg[891]),
    .S(raddr_b_i[0]),
    .X(_2808_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6751_ (.A0(rf_reg[923]),
    .A1(rf_reg[955]),
    .S(raddr_b_i[0]),
    .X(_2809_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6752_ (.Y(_2810_),
    .B1(_2809_),
    .B2(net208),
    .A2(_2808_),
    .A1(net178),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6753_ (.Y(_2811_),
    .A(_2807_),
    .B(_2810_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6754_ (.Y(_2812_),
    .B1(_2811_),
    .B2(net295),
    .A2(_2804_),
    .A1(net300),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6755_ (.B(_2797_),
    .C(_2812_),
    .A(_2788_),
    .Y(rdata_b_o[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6756_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[538]),
    .A1(rf_reg[570]),
    .A2(rf_reg[602]),
    .A3(rf_reg[634]),
    .S1(raddr_b_i[1]),
    .X(_2813_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6757_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[666]),
    .A1(rf_reg[698]),
    .A2(rf_reg[730]),
    .A3(rf_reg[762]),
    .S1(raddr_b_i[1]),
    .X(_2814_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6758_ (.Y(_2815_),
    .B1(_2814_),
    .B2(net218),
    .A2(_2813_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6759_ (.Y(_2816_),
    .A(rf_reg[58]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6760_ (.A0(rf_reg[90]),
    .A1(rf_reg[122]),
    .S(raddr_b_i[0]),
    .X(_2817_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6761_ (.Y(_2818_),
    .A(raddr_b_i[1]),
    .B(_2817_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6762_ (.B1(_2818_),
    .VDD(VDD),
    .Y(_2819_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2816_));
 sg13g2_mux2_1 _6763_ (.A0(rf_reg[154]),
    .A1(rf_reg[186]),
    .S(raddr_b_i[0]),
    .X(_2820_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6764_ (.A0(rf_reg[218]),
    .A1(rf_reg[250]),
    .S(raddr_b_i[0]),
    .X(_2821_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6765_ (.Y(_2822_),
    .B1(_2821_),
    .B2(net186),
    .A2(_2820_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6766_ (.A(net302),
    .B(_2822_),
    .Y(_2823_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6767_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net213),
    .A2(_2819_),
    .Y(_2824_),
    .B1(_2823_));
 sg13g2_mux2_1 _6768_ (.A0(rf_reg[474]),
    .A1(rf_reg[506]),
    .S(raddr_b_i[0]),
    .X(_2825_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6769_ (.A0(rf_reg[346]),
    .A1(rf_reg[378]),
    .S(raddr_b_i[0]),
    .X(_2826_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6770_ (.Y(_2827_),
    .B1(_2826_),
    .B2(net174),
    .A2(_2825_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6771_ (.A0(rf_reg[410]),
    .A1(rf_reg[442]),
    .S(raddr_b_i[0]),
    .X(_2828_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6772_ (.A0(rf_reg[282]),
    .A1(rf_reg[314]),
    .S(raddr_b_i[0]),
    .X(_2829_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6773_ (.Y(_2830_),
    .B1(_2829_),
    .B2(net161),
    .A2(_2828_),
    .A1(net197),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6774_ (.Y(_2831_),
    .A(_2827_),
    .B(_2830_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6775_ (.A0(rf_reg[986]),
    .A1(rf_reg[1018]),
    .S(raddr_b_i[0]),
    .X(_2832_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6776_ (.A0(rf_reg[794]),
    .A1(rf_reg[826]),
    .S(raddr_b_i[0]),
    .X(_2833_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6777_ (.Y(_2834_),
    .B1(_2833_),
    .B2(net161),
    .A2(_2832_),
    .A1(net182),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6778_ (.A0(rf_reg[858]),
    .A1(rf_reg[890]),
    .S(raddr_b_i[0]),
    .X(_2835_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6779_ (.A0(rf_reg[922]),
    .A1(rf_reg[954]),
    .S(raddr_b_i[0]),
    .X(_2836_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6780_ (.Y(_2837_),
    .B1(_2836_),
    .B2(net197),
    .A2(_2835_),
    .A1(net174),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6781_ (.Y(_2838_),
    .A(_2834_),
    .B(_2837_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6782_ (.Y(_2839_),
    .B1(_2838_),
    .B2(net291),
    .A2(_2831_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6783_ (.B(_2824_),
    .C(_2839_),
    .A(_2815_),
    .Y(rdata_b_o[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6784_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[537]),
    .A1(rf_reg[569]),
    .A2(rf_reg[601]),
    .A3(rf_reg[633]),
    .S1(raddr_b_i[1]),
    .X(_2840_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6785_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[665]),
    .A1(rf_reg[697]),
    .A2(rf_reg[729]),
    .A3(rf_reg[761]),
    .S1(raddr_b_i[1]),
    .X(_2841_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6786_ (.Y(_2842_),
    .B1(_2841_),
    .B2(net221),
    .A2(_2840_),
    .A1(net226),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6787_ (.Y(_2843_),
    .A(rf_reg[57]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6788_ (.A0(rf_reg[89]),
    .A1(rf_reg[121]),
    .S(raddr_b_i[0]),
    .X(_2844_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6789_ (.Y(_2845_),
    .A(raddr_b_i[1]),
    .B(_2844_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6790_ (.B1(_2845_),
    .VDD(VDD),
    .Y(_2846_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2843_));
 sg13g2_mux2_1 _6791_ (.A0(rf_reg[153]),
    .A1(rf_reg[185]),
    .S(raddr_b_i[0]),
    .X(_2847_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6792_ (.A0(rf_reg[217]),
    .A1(rf_reg[249]),
    .S(raddr_b_i[0]),
    .X(_2848_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6793_ (.Y(_2849_),
    .B1(_2848_),
    .B2(net188),
    .A2(_2847_),
    .A1(net203),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6794_ (.A(net305),
    .B(_2849_),
    .Y(_2850_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6795_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net216),
    .A2(_2846_),
    .Y(_2851_),
    .B1(_2850_));
 sg13g2_mux2_1 _6796_ (.A0(rf_reg[473]),
    .A1(rf_reg[505]),
    .S(raddr_b_i[0]),
    .X(_2852_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6797_ (.A0(rf_reg[345]),
    .A1(rf_reg[377]),
    .S(raddr_b_i[0]),
    .X(_2853_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6798_ (.Y(_2854_),
    .B1(_2853_),
    .B2(net176),
    .A2(_2852_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6799_ (.A0(rf_reg[409]),
    .A1(rf_reg[441]),
    .S(raddr_b_i[0]),
    .X(_2855_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6800_ (.A0(rf_reg[281]),
    .A1(rf_reg[313]),
    .S(raddr_b_i[0]),
    .X(_2856_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6801_ (.Y(_2857_),
    .B1(_2856_),
    .B2(net163),
    .A2(_2855_),
    .A1(net199),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6802_ (.Y(_2858_),
    .A(_2854_),
    .B(_2857_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6803_ (.A0(rf_reg[985]),
    .A1(rf_reg[1017]),
    .S(raddr_b_i[0]),
    .X(_2859_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6804_ (.A0(rf_reg[793]),
    .A1(rf_reg[825]),
    .S(raddr_b_i[0]),
    .X(_2860_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6805_ (.Y(_2861_),
    .B1(_2860_),
    .B2(net164),
    .A2(_2859_),
    .A1(net184),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6806_ (.A0(rf_reg[857]),
    .A1(rf_reg[889]),
    .S(raddr_b_i[0]),
    .X(_2862_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6807_ (.A0(rf_reg[921]),
    .A1(rf_reg[953]),
    .S(raddr_b_i[0]),
    .X(_2863_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6808_ (.Y(_2864_),
    .B1(_2863_),
    .B2(net200),
    .A2(_2862_),
    .A1(net175),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6809_ (.Y(_2865_),
    .A(_2861_),
    .B(_2864_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6810_ (.Y(_2866_),
    .B1(_2865_),
    .B2(net295),
    .A2(_2858_),
    .A1(net300),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6811_ (.B(_2851_),
    .C(_2866_),
    .A(_2842_),
    .Y(rdata_b_o[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6812_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[536]),
    .A1(rf_reg[568]),
    .A2(rf_reg[600]),
    .A3(rf_reg[632]),
    .S1(raddr_b_i[1]),
    .X(_2867_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6813_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[664]),
    .A1(rf_reg[696]),
    .A2(rf_reg[728]),
    .A3(rf_reg[760]),
    .S1(raddr_b_i[1]),
    .X(_2868_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6814_ (.Y(_2869_),
    .B1(_2868_),
    .B2(net219),
    .A2(_2867_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6815_ (.Y(_2870_),
    .A(rf_reg[56]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6816_ (.A0(rf_reg[88]),
    .A1(rf_reg[120]),
    .S(raddr_b_i[0]),
    .X(_2871_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6817_ (.Y(_2872_),
    .A(raddr_b_i[1]),
    .B(_2871_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6818_ (.B1(_2872_),
    .VDD(VDD),
    .Y(_2873_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2870_));
 sg13g2_mux2_1 _6819_ (.A0(rf_reg[152]),
    .A1(rf_reg[184]),
    .S(raddr_b_i[0]),
    .X(_2874_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6820_ (.A0(rf_reg[216]),
    .A1(rf_reg[248]),
    .S(raddr_b_i[0]),
    .X(_2875_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6821_ (.Y(_2876_),
    .B1(_2875_),
    .B2(net195),
    .A2(_2874_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6822_ (.A(net303),
    .B(_2876_),
    .Y(_2877_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6823_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2873_),
    .Y(_2878_),
    .B1(_2877_));
 sg13g2_mux2_1 _6824_ (.A0(rf_reg[472]),
    .A1(rf_reg[504]),
    .S(raddr_b_i[0]),
    .X(_2879_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6825_ (.A0(rf_reg[344]),
    .A1(rf_reg[376]),
    .S(raddr_b_i[0]),
    .X(_2880_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6826_ (.Y(_2881_),
    .B1(_2880_),
    .B2(net180),
    .A2(_2879_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6827_ (.A0(rf_reg[408]),
    .A1(rf_reg[440]),
    .S(raddr_b_i[0]),
    .X(_2882_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6828_ (.A0(rf_reg[280]),
    .A1(rf_reg[312]),
    .S(raddr_b_i[0]),
    .X(_2883_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6829_ (.Y(_2884_),
    .B1(_2883_),
    .B2(net169),
    .A2(_2882_),
    .A1(net207),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6830_ (.Y(_2885_),
    .A(_2881_),
    .B(_2884_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6831_ (.A0(rf_reg[984]),
    .A1(rf_reg[1016]),
    .S(raddr_b_i[0]),
    .X(_2886_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6832_ (.A0(rf_reg[792]),
    .A1(rf_reg[824]),
    .S(raddr_b_i[0]),
    .X(_2887_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6833_ (.Y(_2888_),
    .B1(_2887_),
    .B2(net168),
    .A2(_2886_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6834_ (.A0(rf_reg[856]),
    .A1(rf_reg[888]),
    .S(raddr_b_i[0]),
    .X(_2889_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6835_ (.A0(rf_reg[920]),
    .A1(rf_reg[952]),
    .S(raddr_b_i[0]),
    .X(_2890_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6836_ (.Y(_2891_),
    .B1(_2890_),
    .B2(net206),
    .A2(_2889_),
    .A1(net179),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6837_ (.Y(_2892_),
    .A(_2888_),
    .B(_2891_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6838_ (.Y(_2893_),
    .B1(_2892_),
    .B2(net293),
    .A2(_2885_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6839_ (.B(_2878_),
    .C(_2893_),
    .A(_2869_),
    .Y(rdata_b_o[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6840_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[535]),
    .A1(rf_reg[567]),
    .A2(rf_reg[599]),
    .A3(rf_reg[631]),
    .S1(raddr_b_i[1]),
    .X(_2894_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6841_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[663]),
    .A1(rf_reg[695]),
    .A2(rf_reg[727]),
    .A3(rf_reg[759]),
    .S1(raddr_b_i[1]),
    .X(_2895_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6842_ (.Y(_2896_),
    .B1(_2895_),
    .B2(net219),
    .A2(_2894_),
    .A1(net224),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6843_ (.Y(_2897_),
    .A(rf_reg[55]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6844_ (.A0(rf_reg[87]),
    .A1(rf_reg[119]),
    .S(raddr_b_i[0]),
    .X(_2898_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6845_ (.Y(_2899_),
    .A(raddr_b_i[1]),
    .B(_2898_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6846_ (.B1(_2899_),
    .VDD(VDD),
    .Y(_2900_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2897_));
 sg13g2_mux2_1 _6847_ (.A0(rf_reg[151]),
    .A1(rf_reg[183]),
    .S(raddr_b_i[0]),
    .X(_2901_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6848_ (.A0(rf_reg[215]),
    .A1(rf_reg[247]),
    .S(raddr_b_i[0]),
    .X(_2902_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6849_ (.Y(_2903_),
    .B1(_2902_),
    .B2(net195),
    .A2(_2901_),
    .A1(net210),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6850_ (.A(net303),
    .B(_2903_),
    .Y(_2904_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6851_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net214),
    .A2(_2900_),
    .Y(_2905_),
    .B1(_2904_));
 sg13g2_mux2_1 _6852_ (.A0(rf_reg[471]),
    .A1(rf_reg[503]),
    .S(raddr_b_i[0]),
    .X(_2906_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6853_ (.A0(rf_reg[343]),
    .A1(rf_reg[375]),
    .S(raddr_b_i[0]),
    .X(_2907_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6854_ (.Y(_2908_),
    .B1(_2907_),
    .B2(net180),
    .A2(_2906_),
    .A1(net191),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6855_ (.A0(rf_reg[407]),
    .A1(rf_reg[439]),
    .S(raddr_b_i[0]),
    .X(_2909_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6856_ (.A0(rf_reg[279]),
    .A1(rf_reg[311]),
    .S(raddr_b_i[0]),
    .X(_2910_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6857_ (.Y(_2911_),
    .B1(_2910_),
    .B2(net168),
    .A2(_2909_),
    .A1(net206),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6858_ (.Y(_2912_),
    .A(_2908_),
    .B(_2911_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6859_ (.A0(rf_reg[983]),
    .A1(rf_reg[1015]),
    .S(raddr_b_i[0]),
    .X(_2913_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6860_ (.A0(rf_reg[791]),
    .A1(rf_reg[823]),
    .S(raddr_b_i[0]),
    .X(_2914_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6861_ (.Y(_2915_),
    .B1(_2914_),
    .B2(net168),
    .A2(_2913_),
    .A1(net192),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6862_ (.A0(rf_reg[855]),
    .A1(rf_reg[887]),
    .S(raddr_b_i[0]),
    .X(_2916_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6863_ (.A0(rf_reg[919]),
    .A1(rf_reg[951]),
    .S(raddr_b_i[0]),
    .X(_2917_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6864_ (.Y(_2918_),
    .B1(_2917_),
    .B2(net208),
    .A2(_2916_),
    .A1(net179),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6865_ (.Y(_2919_),
    .A(_2915_),
    .B(_2918_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6866_ (.Y(_2920_),
    .B1(_2919_),
    .B2(net293),
    .A2(_2912_),
    .A1(net298),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6867_ (.B(_2905_),
    .C(_2920_),
    .A(_2896_),
    .Y(rdata_b_o[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6868_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[534]),
    .A1(rf_reg[566]),
    .A2(rf_reg[598]),
    .A3(rf_reg[630]),
    .S1(raddr_b_i[1]),
    .X(_2921_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux4_1 _6869_ (.S0(raddr_b_i[0]),
    .A0(rf_reg[662]),
    .A1(rf_reg[694]),
    .A2(rf_reg[726]),
    .A3(rf_reg[758]),
    .S1(raddr_b_i[1]),
    .X(_2922_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6870_ (.Y(_2923_),
    .B1(_2922_),
    .B2(net217),
    .A2(_2921_),
    .A1(net222),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6871_ (.Y(_2924_),
    .A(rf_reg[54]),
    .B(raddr_b_i[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6872_ (.A0(rf_reg[86]),
    .A1(rf_reg[118]),
    .S(raddr_b_i[0]),
    .X(_2925_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6873_ (.Y(_2926_),
    .A(raddr_b_i[1]),
    .B(_2925_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _6874_ (.B1(_2926_),
    .VDD(VDD),
    .Y(_2927_),
    .VSS(VSS),
    .A1(raddr_b_i[1]),
    .A2(_2924_));
 sg13g2_mux2_1 _6875_ (.A0(rf_reg[150]),
    .A1(rf_reg[182]),
    .S(raddr_b_i[0]),
    .X(_2928_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6876_ (.A0(rf_reg[214]),
    .A1(rf_reg[246]),
    .S(raddr_b_i[0]),
    .X(_2929_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6877_ (.Y(_2930_),
    .B1(_2929_),
    .B2(net186),
    .A2(_2928_),
    .A1(net202),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6878_ (.A(net301),
    .B(_2930_),
    .Y(_2931_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _6879_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net212),
    .A2(_2927_),
    .Y(_2932_),
    .B1(_2931_));
 sg13g2_mux2_1 _6880_ (.A0(rf_reg[470]),
    .A1(rf_reg[502]),
    .S(raddr_b_i[0]),
    .X(_2933_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6881_ (.A0(rf_reg[342]),
    .A1(rf_reg[374]),
    .S(raddr_b_i[0]),
    .X(_2934_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6882_ (.Y(_2935_),
    .B1(_2934_),
    .B2(net173),
    .A2(_2933_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6883_ (.A0(rf_reg[406]),
    .A1(rf_reg[438]),
    .S(raddr_b_i[0]),
    .X(_2936_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6884_ (.A0(rf_reg[278]),
    .A1(rf_reg[310]),
    .S(raddr_b_i[0]),
    .X(_2937_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6885_ (.Y(_2938_),
    .B1(_2937_),
    .B2(net162),
    .A2(_2936_),
    .A1(net198),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6886_ (.Y(_2939_),
    .A(_2935_),
    .B(_2938_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6887_ (.A0(rf_reg[982]),
    .A1(rf_reg[1014]),
    .S(raddr_b_i[0]),
    .X(_2940_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6888_ (.A0(rf_reg[790]),
    .A1(rf_reg[822]),
    .S(raddr_b_i[0]),
    .X(_2941_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6889_ (.Y(_2942_),
    .B1(_2941_),
    .B2(net162),
    .A2(_2940_),
    .A1(net183),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6890_ (.A0(rf_reg[854]),
    .A1(rf_reg[886]),
    .S(raddr_b_i[0]),
    .X(_2943_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6891_ (.A0(rf_reg[918]),
    .A1(rf_reg[950]),
    .S(raddr_b_i[0]),
    .X(_2944_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6892_ (.Y(_2945_),
    .B1(_2944_),
    .B2(net198),
    .A2(_2943_),
    .A1(net173),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _6893_ (.Y(_2946_),
    .A(_2942_),
    .B(_2945_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _6894_ (.Y(_2947_),
    .B1(_2946_),
    .B2(net291),
    .A2(_2939_),
    .A1(net296),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _6895_ (.B(_2932_),
    .C(_2947_),
    .A(_2923_),
    .Y(rdata_b_o[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(net115),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 _6897_ (.Y(_2949_),
    .A(waddr_a_i[0]),
    .B(waddr_a_i[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _6898_ (.B(we_a_i),
    .C(waddr_a_i[2]),
    .A(waddr_a_i[4]),
    .Y(_2950_),
    .VDD(VDD),
    .VSS(VSS),
    .D(waddr_a_i[1]));
 sg13g2_nor2_2 _6899_ (.A(_2949_),
    .B(_2950_),
    .Y(_2951_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(net115),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6901_ (.A0(rf_reg[1000]),
    .A1(net341),
    .S(net156),
    .X(_0000_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_3161_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6903_ (.A0(rf_reg[1001]),
    .A1(net347),
    .S(net156),
    .X(_0001_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(net110),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6905_ (.A0(rf_reg[1002]),
    .A1(net327),
    .S(net158),
    .X(_0002_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net109),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6907_ (.A0(rf_reg[1003]),
    .A1(net317),
    .S(net160),
    .X(_0003_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net110),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6909_ (.A0(rf_reg[1004]),
    .A1(net322),
    .S(net156),
    .X(_0004_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net110),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6911_ (.A0(rf_reg[1005]),
    .A1(net345),
    .S(net159),
    .X(_0005_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout105 (.A(_3166_),
    .X(net105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6913_ (.A0(rf_reg[1006]),
    .A1(net321),
    .S(net158),
    .X(_0006_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6915_ (.A0(rf_reg[1007]),
    .A1(net332),
    .S(net158),
    .X(_0007_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net104),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6917_ (.A0(rf_reg[1008]),
    .A1(net320),
    .S(net159),
    .X(_0008_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6919_ (.A0(rf_reg[1009]),
    .A1(net330),
    .S(net157),
    .X(_0009_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net102),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 _6921_ (.Y(_2963_),
    .B(waddr_a_i[0]),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(waddr_a_i[3]));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(_3171_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 _6923_ (.A(waddr_a_i[4]),
    .B_N(we_a_i),
    .Y(_2965_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _6924_ (.A(waddr_a_i[2]),
    .B_N(waddr_a_i[1]),
    .Y(_2966_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 _6925_ (.Y(_2967_),
    .A(_2965_),
    .B(_2966_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _6926_ (.A(_2963_),
    .B(_2967_),
    .Y(_2968_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net100),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6928_ (.A0(rf_reg[100]),
    .A1(net337),
    .S(net61),
    .X(_0010_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(net99),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(net100),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6931_ (.A0(rf_reg[1010]),
    .A1(net318),
    .S(net160),
    .X(_0011_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net97),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6933_ (.A0(rf_reg[1011]),
    .A1(net325),
    .S(net160),
    .X(_0012_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout95 (.A(_3176_),
    .X(net95),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6935_ (.A0(rf_reg[1012]),
    .A1(net344),
    .S(net159),
    .X(_0013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(net95),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6937_ (.A0(rf_reg[1013]),
    .A1(net334),
    .S(net157),
    .X(_0014_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net94),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6939_ (.A0(rf_reg[1014]),
    .A1(net338),
    .S(net157),
    .X(_0015_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net95),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6941_ (.A0(rf_reg[1015]),
    .A1(net324),
    .S(net160),
    .X(_0016_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net92),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6943_ (.A0(rf_reg[1016]),
    .A1(net336),
    .S(net159),
    .X(_0017_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout90 (.A(_3181_),
    .X(net90),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6945_ (.A0(rf_reg[1017]),
    .A1(net333),
    .S(net158),
    .X(_0018_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net90),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6947_ (.A0(rf_reg[1018]),
    .A1(net343),
    .S(net156),
    .X(_0019_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(net89),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6949_ (.A0(rf_reg[1019]),
    .A1(net316),
    .S(net159),
    .X(_0020_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(net90),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6951_ (.A0(rf_reg[101]),
    .A1(net342),
    .S(net63),
    .X(_0021_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(net87),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout85 (.A(_3185_),
    .X(net85),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6954_ (.A0(rf_reg[1020]),
    .A1(net339),
    .S(net159),
    .X(_0022_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net85),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6956_ (.A0(rf_reg[1021]),
    .A1(net335),
    .S(net156),
    .X(_0023_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(net84),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6958_ (.A0(rf_reg[1022]),
    .A1(net319),
    .S(net157),
    .X(_0024_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(net85),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6960_ (.A0(rf_reg[1023]),
    .A1(net323),
    .S(net156),
    .X(_0025_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(net82),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6962_ (.A0(rf_reg[102]),
    .A1(net326),
    .S(net61),
    .X(_0026_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout80 (.A(_3189_),
    .X(net80),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6964_ (.A0(rf_reg[103]),
    .A1(net340),
    .S(net63),
    .X(_0027_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(net80),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6966_ (.A0(rf_reg[104]),
    .A1(net341),
    .S(net61),
    .X(_0028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(net79),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6968_ (.A0(rf_reg[105]),
    .A1(net347),
    .S(net61),
    .X(_0029_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(net80),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6970_ (.A0(rf_reg[106]),
    .A1(net327),
    .S(net62),
    .X(_0030_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(net77),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6972_ (.A0(rf_reg[107]),
    .A1(net317),
    .S(net64),
    .X(_0031_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_3193_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6974_ (.A0(rf_reg[108]),
    .A1(net322),
    .S(net62),
    .X(_0032_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(net75),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6976_ (.A0(rf_reg[109]),
    .A1(net345),
    .S(net63),
    .X(_0033_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_3193_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6979_ (.A0(rf_reg[110]),
    .A1(net321),
    .S(net64),
    .X(_0034_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(net73),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6981_ (.A0(rf_reg[111]),
    .A1(net332),
    .S(net64),
    .X(_0035_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout70 (.A(_1048_),
    .X(net70),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6983_ (.A0(rf_reg[112]),
    .A1(net320),
    .S(net63),
    .X(_0036_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(net70),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6985_ (.A0(rf_reg[113]),
    .A1(net330),
    .S(net61),
    .X(_0037_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(net69),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6987_ (.A0(rf_reg[114]),
    .A1(net318),
    .S(net64),
    .X(_0038_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(net70),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6989_ (.A0(rf_reg[115]),
    .A1(net325),
    .S(net64),
    .X(_0039_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(net67),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6991_ (.A0(rf_reg[116]),
    .A1(net344),
    .S(net63),
    .X(_0040_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout65 (.A(_2968_),
    .X(net65),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6993_ (.A0(rf_reg[117]),
    .A1(net334),
    .S(net61),
    .X(_0041_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(net65),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6995_ (.A0(rf_reg[118]),
    .A1(net338),
    .S(net61),
    .X(_0042_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net64),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _6997_ (.A0(rf_reg[119]),
    .A1(net324),
    .S(net63),
    .X(_0043_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net65),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net62),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7000_ (.A0(rf_reg[120]),
    .A1(net336),
    .S(net65),
    .X(_0044_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout60 (.A(_3020_),
    .X(net60),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7002_ (.A0(rf_reg[121]),
    .A1(net333),
    .S(net62),
    .X(_0045_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(net60),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7004_ (.A0(rf_reg[122]),
    .A1(net343),
    .S(net62),
    .X(_0046_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(net60),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7006_ (.A0(rf_reg[123]),
    .A1(net316),
    .S(net65),
    .X(_0047_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(net60),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7008_ (.A0(rf_reg[124]),
    .A1(net339),
    .S(net63),
    .X(_0048_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7010_ (.A0(rf_reg[125]),
    .A1(net335),
    .S(net62),
    .X(_0049_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(_3028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7012_ (.A0(rf_reg[126]),
    .A1(net319),
    .S(net62),
    .X(_0050_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7014_ (.A0(rf_reg[127]),
    .A1(net323),
    .S(net62),
    .X(_0051_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 _7016_ (.VSS(VSS),
    .VDD(VDD),
    .X(_3016_),
    .B(waddr_a_i[3]),
    .A(waddr_a_i[0]));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _7018_ (.A(waddr_a_i[1]),
    .B_N(waddr_a_i[2]),
    .Y(_3018_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 _7019_ (.Y(_3019_),
    .A(_2965_),
    .B(_3018_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _7020_ (.VSS(VSS),
    .VDD(VDD),
    .X(_3020_),
    .B(_3019_),
    .A(_3016_));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(net52),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout50 (.A(_3038_),
    .X(net50),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7023_ (.A0(net328),
    .A1(rf_reg[128]),
    .S(net58),
    .X(_0052_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(net50),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7025_ (.A0(net329),
    .A1(rf_reg[129]),
    .S(net58),
    .X(_0053_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(net50),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7027_ (.A0(net346),
    .A1(rf_reg[130]),
    .S(net57),
    .X(_0054_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(net50),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7029_ (.A0(net331),
    .A1(rf_reg[131]),
    .S(net59),
    .X(_0055_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7030_ (.A0(net337),
    .A1(rf_reg[132]),
    .S(net56),
    .X(_0056_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7031_ (.A0(net342),
    .A1(rf_reg[133]),
    .S(net59),
    .X(_0057_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7032_ (.A0(net326),
    .A1(rf_reg[134]),
    .S(net56),
    .X(_0058_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7033_ (.A0(net340),
    .A1(rf_reg[135]),
    .S(net59),
    .X(_0059_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7034_ (.A0(net341),
    .A1(rf_reg[136]),
    .S(net56),
    .X(_0060_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7035_ (.A0(net347),
    .A1(rf_reg[137]),
    .S(net56),
    .X(_0061_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(net47),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7037_ (.A0(net327),
    .A1(rf_reg[138]),
    .S(net57),
    .X(_0062_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7038_ (.A0(net317),
    .A1(rf_reg[139]),
    .S(net58),
    .X(_0063_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7039_ (.A0(net322),
    .A1(rf_reg[140]),
    .S(net57),
    .X(_0064_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7040_ (.A0(net345),
    .A1(rf_reg[141]),
    .S(net59),
    .X(_0065_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7041_ (.A0(net321),
    .A1(rf_reg[142]),
    .S(net58),
    .X(_0066_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7042_ (.A0(net332),
    .A1(rf_reg[143]),
    .S(net58),
    .X(_0067_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7043_ (.A0(net320),
    .A1(rf_reg[144]),
    .S(net58),
    .X(_0068_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7044_ (.A0(net330),
    .A1(rf_reg[145]),
    .S(net56),
    .X(_0069_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7045_ (.A0(net318),
    .A1(rf_reg[146]),
    .S(net57),
    .X(_0070_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7046_ (.A0(net325),
    .A1(rf_reg[147]),
    .S(net58),
    .X(_0071_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout45 (.X(net45),
    .A(_3045_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7048_ (.A0(net344),
    .A1(rf_reg[148]),
    .S(net59),
    .X(_0072_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7049_ (.A0(net334),
    .A1(rf_reg[149]),
    .S(net56),
    .X(_0073_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7050_ (.A0(net338),
    .A1(rf_reg[150]),
    .S(net56),
    .X(_0074_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7051_ (.A0(net324),
    .A1(rf_reg[151]),
    .S(net59),
    .X(_0075_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7052_ (.A0(net336),
    .A1(rf_reg[152]),
    .S(net59),
    .X(_0076_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7053_ (.A0(net333),
    .A1(rf_reg[153]),
    .S(net60),
    .X(_0077_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7054_ (.A0(net343),
    .A1(rf_reg[154]),
    .S(net57),
    .X(_0078_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7055_ (.A0(net316),
    .A1(rf_reg[155]),
    .S(net58),
    .X(_0079_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7056_ (.A0(net339),
    .A1(rf_reg[156]),
    .S(net59),
    .X(_0080_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7057_ (.A0(net335),
    .A1(rf_reg[157]),
    .S(net56),
    .X(_0081_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7058_ (.A0(net319),
    .A1(rf_reg[158]),
    .S(net57),
    .X(_0082_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7059_ (.A0(net323),
    .A1(rf_reg[159]),
    .S(net57),
    .X(_0083_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7060_ (.A(_2963_),
    .B(_3019_),
    .Y(_3028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(net45),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7062_ (.A0(rf_reg[160]),
    .A1(net328),
    .S(net53),
    .X(_0084_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7063_ (.A0(rf_reg[161]),
    .A1(net329),
    .S(net53),
    .X(_0085_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7064_ (.A0(rf_reg[162]),
    .A1(net346),
    .S(net52),
    .X(_0086_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7065_ (.A0(rf_reg[163]),
    .A1(net331),
    .S(net54),
    .X(_0087_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(net44),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7067_ (.A0(rf_reg[164]),
    .A1(net337),
    .S(net51),
    .X(_0088_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net45),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7069_ (.A0(rf_reg[165]),
    .A1(net342),
    .S(net53),
    .X(_0089_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(net45),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7071_ (.A0(rf_reg[166]),
    .A1(net326),
    .S(net51),
    .X(_0090_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_3053_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7073_ (.A0(rf_reg[167]),
    .A1(net340),
    .S(net53),
    .X(_0091_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7074_ (.A0(rf_reg[168]),
    .A1(net341),
    .S(net51),
    .X(_0092_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7075_ (.A0(rf_reg[169]),
    .A1(net347),
    .S(net51),
    .X(_0093_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(net40),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7077_ (.A0(rf_reg[170]),
    .A1(net327),
    .S(net55),
    .X(_0094_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7078_ (.A0(rf_reg[171]),
    .A1(net317),
    .S(net53),
    .X(_0095_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7079_ (.A0(rf_reg[172]),
    .A1(net322),
    .S(net55),
    .X(_0096_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7080_ (.A0(rf_reg[173]),
    .A1(net345),
    .S(net54),
    .X(_0097_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7081_ (.A0(rf_reg[174]),
    .A1(net321),
    .S(net52),
    .X(_0098_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7082_ (.A0(rf_reg[175]),
    .A1(net332),
    .S(net52),
    .X(_0099_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7083_ (.A0(rf_reg[176]),
    .A1(net320),
    .S(net53),
    .X(_0100_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7084_ (.A0(rf_reg[177]),
    .A1(net330),
    .S(net51),
    .X(_0101_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7085_ (.A0(rf_reg[178]),
    .A1(net318),
    .S(net52),
    .X(_0102_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7086_ (.A0(rf_reg[179]),
    .A1(net325),
    .S(net53),
    .X(_0103_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(net40),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7088_ (.A0(rf_reg[180]),
    .A1(net344),
    .S(net54),
    .X(_0104_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7089_ (.A0(rf_reg[181]),
    .A1(net334),
    .S(net51),
    .X(_0105_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7090_ (.A0(rf_reg[182]),
    .A1(net338),
    .S(net51),
    .X(_0106_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7091_ (.A0(rf_reg[183]),
    .A1(net324),
    .S(net54),
    .X(_0107_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7092_ (.A0(rf_reg[184]),
    .A1(net336),
    .S(net54),
    .X(_0108_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7093_ (.A0(rf_reg[185]),
    .A1(net333),
    .S(net55),
    .X(_0109_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7094_ (.A0(rf_reg[186]),
    .A1(net343),
    .S(net52),
    .X(_0110_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7095_ (.A0(rf_reg[187]),
    .A1(net316),
    .S(net53),
    .X(_0111_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7096_ (.A0(rf_reg[188]),
    .A1(net339),
    .S(net54),
    .X(_0112_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7097_ (.A0(rf_reg[189]),
    .A1(net335),
    .S(net51),
    .X(_0113_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7098_ (.A0(rf_reg[190]),
    .A1(net319),
    .S(net52),
    .X(_0114_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7099_ (.A0(rf_reg[191]),
    .A1(net323),
    .S(net52),
    .X(_0115_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(net40),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _7101_ (.B(waddr_a_i[1]),
    .C(_2965_),
    .A(waddr_a_i[2]),
    .Y(_3037_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7102_ (.A(_3016_),
    .B(_3037_),
    .Y(_3038_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout36 (.X(net36),
    .A(net40),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7104_ (.A0(rf_reg[192]),
    .A1(net328),
    .S(net49),
    .X(_0116_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(_3058_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7106_ (.A0(rf_reg[193]),
    .A1(net329),
    .S(net49),
    .X(_0117_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7108_ (.A0(rf_reg[194]),
    .A1(net346),
    .S(net46),
    .X(_0118_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7110_ (.A0(rf_reg[195]),
    .A1(net331),
    .S(net48),
    .X(_0119_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7111_ (.A0(rf_reg[196]),
    .A1(net337),
    .S(net46),
    .X(_0120_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7112_ (.A0(rf_reg[197]),
    .A1(net342),
    .S(net48),
    .X(_0121_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7113_ (.A0(rf_reg[198]),
    .A1(net326),
    .S(net47),
    .X(_0122_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7114_ (.A0(rf_reg[199]),
    .A1(net340),
    .S(net48),
    .X(_0123_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7115_ (.A0(rf_reg[200]),
    .A1(net341),
    .S(net46),
    .X(_0124_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7116_ (.A0(rf_reg[201]),
    .A1(net347),
    .S(net46),
    .X(_0125_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout32 (.X(net32),
    .A(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7118_ (.A0(rf_reg[202]),
    .A1(net327),
    .S(net47),
    .X(_0126_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7119_ (.A0(rf_reg[203]),
    .A1(net317),
    .S(net49),
    .X(_0127_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7120_ (.A0(rf_reg[204]),
    .A1(net322),
    .S(net47),
    .X(_0128_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7121_ (.A0(rf_reg[205]),
    .A1(net345),
    .S(net48),
    .X(_0129_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7122_ (.A0(rf_reg[206]),
    .A1(net321),
    .S(net49),
    .X(_0130_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7123_ (.A0(rf_reg[207]),
    .A1(net332),
    .S(net49),
    .X(_0131_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7124_ (.A0(rf_reg[208]),
    .A1(net320),
    .S(net48),
    .X(_0132_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7125_ (.A0(rf_reg[209]),
    .A1(net330),
    .S(net46),
    .X(_0133_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7126_ (.A0(rf_reg[210]),
    .A1(net318),
    .S(net49),
    .X(_0134_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7127_ (.A0(rf_reg[211]),
    .A1(net325),
    .S(net49),
    .X(_0135_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout31 (.X(net31),
    .A(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7129_ (.A0(rf_reg[212]),
    .A1(net344),
    .S(net50),
    .X(_0136_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7130_ (.A0(rf_reg[213]),
    .A1(net334),
    .S(net46),
    .X(_0137_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7131_ (.A0(rf_reg[214]),
    .A1(net338),
    .S(net46),
    .X(_0138_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7132_ (.A0(rf_reg[215]),
    .A1(net324),
    .S(net48),
    .X(_0139_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7133_ (.A0(rf_reg[216]),
    .A1(net336),
    .S(net48),
    .X(_0140_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7134_ (.A0(rf_reg[217]),
    .A1(net333),
    .S(net47),
    .X(_0141_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7135_ (.A0(rf_reg[218]),
    .A1(net343),
    .S(net47),
    .X(_0142_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7136_ (.A0(rf_reg[219]),
    .A1(net316),
    .S(net49),
    .X(_0143_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7137_ (.A0(rf_reg[220]),
    .A1(net339),
    .S(net48),
    .X(_0144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7138_ (.A0(rf_reg[221]),
    .A1(net335),
    .S(net46),
    .X(_0145_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7139_ (.A0(rf_reg[222]),
    .A1(net319),
    .S(net47),
    .X(_0146_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7140_ (.A0(rf_reg[223]),
    .A1(net323),
    .S(net47),
    .X(_0147_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7141_ (.A(_2963_),
    .B(_3037_),
    .Y(_3045_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout30 (.X(net30),
    .A(_3063_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7143_ (.A0(rf_reg[224]),
    .A1(net328),
    .S(net43),
    .X(_0148_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7144_ (.A0(rf_reg[225]),
    .A1(net329),
    .S(net43),
    .X(_0149_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7145_ (.A0(rf_reg[226]),
    .A1(net346),
    .S(net41),
    .X(_0150_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7146_ (.A0(rf_reg[227]),
    .A1(net331),
    .S(net44),
    .X(_0151_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7147_ (.A0(rf_reg[228]),
    .A1(net337),
    .S(net41),
    .X(_0152_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7148_ (.A0(rf_reg[229]),
    .A1(net342),
    .S(net44),
    .X(_0153_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7149_ (.A0(rf_reg[230]),
    .A1(net326),
    .S(net42),
    .X(_0154_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7150_ (.A0(rf_reg[231]),
    .A1(net340),
    .S(net44),
    .X(_0155_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7151_ (.A0(rf_reg[232]),
    .A1(net341),
    .S(net41),
    .X(_0156_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7152_ (.A0(rf_reg[233]),
    .A1(net347),
    .S(net41),
    .X(_0157_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 fanout29 (.A(net30),
    .X(net29),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7154_ (.A0(rf_reg[234]),
    .A1(net327),
    .S(net42),
    .X(_0158_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7155_ (.A0(rf_reg[235]),
    .A1(net317),
    .S(net43),
    .X(_0159_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7156_ (.A0(rf_reg[236]),
    .A1(net322),
    .S(net42),
    .X(_0160_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7157_ (.A0(rf_reg[237]),
    .A1(net345),
    .S(net44),
    .X(_0161_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7158_ (.A0(rf_reg[238]),
    .A1(net321),
    .S(net43),
    .X(_0162_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7159_ (.A0(rf_reg[239]),
    .A1(net332),
    .S(net43),
    .X(_0163_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7160_ (.A0(rf_reg[240]),
    .A1(net320),
    .S(net43),
    .X(_0164_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7161_ (.A0(rf_reg[241]),
    .A1(net330),
    .S(net41),
    .X(_0165_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7162_ (.A0(rf_reg[242]),
    .A1(net318),
    .S(net43),
    .X(_0166_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7163_ (.A0(rf_reg[243]),
    .A1(net325),
    .S(net43),
    .X(_0167_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout28 (.X(net28),
    .A(net29),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7165_ (.A0(rf_reg[244]),
    .A1(net344),
    .S(net45),
    .X(_0168_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7166_ (.A0(rf_reg[245]),
    .A1(net334),
    .S(net41),
    .X(_0169_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7167_ (.A0(rf_reg[246]),
    .A1(net338),
    .S(net41),
    .X(_0170_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7168_ (.A0(rf_reg[247]),
    .A1(net324),
    .S(net45),
    .X(_0171_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7169_ (.A0(rf_reg[248]),
    .A1(net336),
    .S(net44),
    .X(_0172_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7170_ (.A0(rf_reg[249]),
    .A1(net333),
    .S(net42),
    .X(_0173_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7171_ (.A0(rf_reg[250]),
    .A1(net343),
    .S(net42),
    .X(_0174_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7172_ (.A0(rf_reg[251]),
    .A1(net316),
    .S(net44),
    .X(_0175_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7173_ (.A0(rf_reg[252]),
    .A1(net339),
    .S(net44),
    .X(_0176_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7174_ (.A0(rf_reg[253]),
    .A1(net335),
    .S(net41),
    .X(_0177_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7175_ (.A0(rf_reg[254]),
    .A1(net319),
    .S(net42),
    .X(_0178_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7176_ (.A0(rf_reg[255]),
    .A1(net323),
    .S(net42),
    .X(_0179_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_2 _7177_ (.Y(_3049_),
    .B(waddr_a_i[3]),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(waddr_a_i[0]));
 sg13g2_buf_4 fanout27 (.X(net27),
    .A(net30),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7179_ (.A(waddr_a_i[2]),
    .B(waddr_a_i[1]),
    .Y(_3051_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _7180_ (.A(_2965_),
    .B(_3051_),
    .X(_3052_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _7181_ (.Y(_3053_),
    .B(_3052_),
    .A_N(_3049_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(net30),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout25 (.A(_3065_),
    .X(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7184_ (.A0(net328),
    .A1(rf_reg[256]),
    .S(net39),
    .X(_0180_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7185_ (.A0(net329),
    .A1(rf_reg[257]),
    .S(net39),
    .X(_0181_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7186_ (.A0(net346),
    .A1(rf_reg[258]),
    .S(net36),
    .X(_0182_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7187_ (.A0(net331),
    .A1(rf_reg[259]),
    .S(net38),
    .X(_0183_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7188_ (.A0(net337),
    .A1(rf_reg[260]),
    .S(net36),
    .X(_0184_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7189_ (.A0(net342),
    .A1(rf_reg[261]),
    .S(net38),
    .X(_0185_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7190_ (.A0(net326),
    .A1(rf_reg[262]),
    .S(net37),
    .X(_0186_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7191_ (.A0(net340),
    .A1(rf_reg[263]),
    .S(net38),
    .X(_0187_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7192_ (.A0(net341),
    .A1(rf_reg[264]),
    .S(net37),
    .X(_0188_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7193_ (.A0(net347),
    .A1(rf_reg[265]),
    .S(net36),
    .X(_0189_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout24 (.X(net24),
    .A(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7195_ (.A0(net327),
    .A1(rf_reg[266]),
    .S(net37),
    .X(_0190_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7196_ (.A0(net317),
    .A1(rf_reg[267]),
    .S(net39),
    .X(_0191_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7197_ (.A0(net322),
    .A1(rf_reg[268]),
    .S(net37),
    .X(_0192_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7198_ (.A0(net345),
    .A1(rf_reg[269]),
    .S(net38),
    .X(_0193_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7199_ (.A0(net321),
    .A1(rf_reg[270]),
    .S(net39),
    .X(_0194_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7200_ (.A0(net332),
    .A1(rf_reg[271]),
    .S(net39),
    .X(_0195_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7201_ (.A0(net320),
    .A1(rf_reg[272]),
    .S(net39),
    .X(_0196_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7202_ (.A0(net330),
    .A1(rf_reg[273]),
    .S(net36),
    .X(_0197_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7203_ (.A0(net318),
    .A1(rf_reg[274]),
    .S(net39),
    .X(_0198_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7204_ (.A0(net325),
    .A1(rf_reg[275]),
    .S(net39),
    .X(_0199_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(net24),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7206_ (.A0(net344),
    .A1(rf_reg[276]),
    .S(net38),
    .X(_0200_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7207_ (.A0(net334),
    .A1(rf_reg[277]),
    .S(net36),
    .X(_0201_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7208_ (.A0(net338),
    .A1(rf_reg[278]),
    .S(net36),
    .X(_0202_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7209_ (.A0(net324),
    .A1(rf_reg[279]),
    .S(net40),
    .X(_0203_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7210_ (.A0(net336),
    .A1(rf_reg[280]),
    .S(net38),
    .X(_0204_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7211_ (.A0(net333),
    .A1(rf_reg[281]),
    .S(net37),
    .X(_0205_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7212_ (.A0(net343),
    .A1(rf_reg[282]),
    .S(net36),
    .X(_0206_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7213_ (.A0(net316),
    .A1(rf_reg[283]),
    .S(net38),
    .X(_0207_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7214_ (.A0(net339),
    .A1(rf_reg[284]),
    .S(net38),
    .X(_0208_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7215_ (.A0(net335),
    .A1(rf_reg[285]),
    .S(net36),
    .X(_0209_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7216_ (.A0(net319),
    .A1(rf_reg[286]),
    .S(net37),
    .X(_0210_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7217_ (.A0(net323),
    .A1(rf_reg[287]),
    .S(net37),
    .X(_0211_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _7218_ (.Y(_3058_),
    .B(_3052_),
    .A_N(_2949_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout22 (.X(net22),
    .A(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout21 (.X(net21),
    .A(net22),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7221_ (.A0(net328),
    .A1(rf_reg[288]),
    .S(net34),
    .X(_0212_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7222_ (.A0(net329),
    .A1(rf_reg[289]),
    .S(net34),
    .X(_0213_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7223_ (.A0(net346),
    .A1(rf_reg[290]),
    .S(net31),
    .X(_0214_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7224_ (.A0(net331),
    .A1(rf_reg[291]),
    .S(net33),
    .X(_0215_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7225_ (.A0(net337),
    .A1(rf_reg[292]),
    .S(net31),
    .X(_0216_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7226_ (.A0(net342),
    .A1(rf_reg[293]),
    .S(net33),
    .X(_0217_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7227_ (.A0(net326),
    .A1(rf_reg[294]),
    .S(net32),
    .X(_0218_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7228_ (.A0(net340),
    .A1(rf_reg[295]),
    .S(net33),
    .X(_0219_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7229_ (.A0(net341),
    .A1(rf_reg[296]),
    .S(net32),
    .X(_0220_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7230_ (.A0(net347),
    .A1(rf_reg[297]),
    .S(net31),
    .X(_0221_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout20 (.X(net20),
    .A(_3070_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7232_ (.A0(net327),
    .A1(rf_reg[298]),
    .S(net32),
    .X(_0222_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7233_ (.A0(net317),
    .A1(rf_reg[299]),
    .S(net34),
    .X(_0223_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7234_ (.A0(net322),
    .A1(rf_reg[300]),
    .S(net32),
    .X(_0224_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7235_ (.A0(net345),
    .A1(rf_reg[301]),
    .S(net33),
    .X(_0225_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7236_ (.A0(net321),
    .A1(rf_reg[302]),
    .S(net34),
    .X(_0226_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7237_ (.A0(net332),
    .A1(rf_reg[303]),
    .S(net34),
    .X(_0227_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7238_ (.A0(net320),
    .A1(rf_reg[304]),
    .S(net33),
    .X(_0228_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7239_ (.A0(net330),
    .A1(rf_reg[305]),
    .S(net31),
    .X(_0229_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7240_ (.A0(net318),
    .A1(rf_reg[306]),
    .S(net34),
    .X(_0230_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7241_ (.A0(net325),
    .A1(rf_reg[307]),
    .S(net34),
    .X(_0231_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout19 (.X(net19),
    .A(net20),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7243_ (.A0(net344),
    .A1(rf_reg[308]),
    .S(net33),
    .X(_0232_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7244_ (.A0(net334),
    .A1(rf_reg[309]),
    .S(net31),
    .X(_0233_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7245_ (.A0(net338),
    .A1(rf_reg[310]),
    .S(net31),
    .X(_0234_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7246_ (.A0(net324),
    .A1(rf_reg[311]),
    .S(net35),
    .X(_0235_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7247_ (.A0(net336),
    .A1(rf_reg[312]),
    .S(net33),
    .X(_0236_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7248_ (.A0(net333),
    .A1(rf_reg[313]),
    .S(net32),
    .X(_0237_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7249_ (.A0(net343),
    .A1(rf_reg[314]),
    .S(net31),
    .X(_0238_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7250_ (.A0(net316),
    .A1(rf_reg[315]),
    .S(net35),
    .X(_0239_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7251_ (.A0(net339),
    .A1(rf_reg[316]),
    .S(net33),
    .X(_0240_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7252_ (.A0(net335),
    .A1(rf_reg[317]),
    .S(net31),
    .X(_0241_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7253_ (.A0(net319),
    .A1(rf_reg[318]),
    .S(net32),
    .X(_0242_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7254_ (.A0(net323),
    .A1(rf_reg[319]),
    .S(net32),
    .X(_0243_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7255_ (.A(_2967_),
    .B(_3049_),
    .Y(_3063_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout18 (.X(net18),
    .A(net19),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7257_ (.A0(rf_reg[320]),
    .A1(net328),
    .S(net29),
    .X(_0244_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7258_ (.A0(rf_reg[321]),
    .A1(net329),
    .S(net29),
    .X(_0245_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7259_ (.A0(rf_reg[322]),
    .A1(net346),
    .S(net26),
    .X(_0246_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7260_ (.A0(rf_reg[323]),
    .A1(net331),
    .S(net28),
    .X(_0247_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7261_ (.A0(rf_reg[324]),
    .A1(net337),
    .S(net26),
    .X(_0248_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7262_ (.A0(rf_reg[325]),
    .A1(net342),
    .S(net28),
    .X(_0249_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7263_ (.A0(rf_reg[326]),
    .A1(net326),
    .S(net27),
    .X(_0250_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7264_ (.A0(rf_reg[327]),
    .A1(net340),
    .S(net28),
    .X(_0251_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7265_ (.A0(rf_reg[328]),
    .A1(net341),
    .S(net27),
    .X(_0252_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7266_ (.A0(rf_reg[329]),
    .A1(net347),
    .S(net26),
    .X(_0253_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _7267_ (.Y(_3065_),
    .B(_3052_),
    .A_N(_2963_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout17 (.X(net17),
    .A(net20),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout16 (.X(net16),
    .A(net20),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7270_ (.A0(net328),
    .A1(rf_reg[32]),
    .S(net24),
    .X(_0254_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout15 (.X(net15),
    .A(_3074_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7272_ (.A0(rf_reg[330]),
    .A1(net327),
    .S(net27),
    .X(_0255_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7273_ (.A0(rf_reg[331]),
    .A1(net317),
    .S(net29),
    .X(_0256_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7274_ (.A0(rf_reg[332]),
    .A1(net322),
    .S(net27),
    .X(_0257_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7275_ (.A0(rf_reg[333]),
    .A1(net345),
    .S(net28),
    .X(_0258_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7276_ (.A0(rf_reg[334]),
    .A1(net321),
    .S(net27),
    .X(_0259_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7277_ (.A0(rf_reg[335]),
    .A1(net332),
    .S(net29),
    .X(_0260_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7278_ (.A0(rf_reg[336]),
    .A1(net320),
    .S(net29),
    .X(_0261_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7279_ (.A0(rf_reg[337]),
    .A1(net330),
    .S(net26),
    .X(_0262_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7280_ (.A0(rf_reg[338]),
    .A1(net318),
    .S(net29),
    .X(_0263_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7281_ (.A0(rf_reg[339]),
    .A1(net325),
    .S(net29),
    .X(_0264_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7282_ (.A0(net329),
    .A1(rf_reg[33]),
    .S(net24),
    .X(_0265_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout14 (.X(net14),
    .A(net15),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7284_ (.A0(rf_reg[340]),
    .A1(net344),
    .S(net28),
    .X(_0266_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7285_ (.A0(rf_reg[341]),
    .A1(net334),
    .S(net26),
    .X(_0267_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7286_ (.A0(rf_reg[342]),
    .A1(net338),
    .S(net26),
    .X(_0268_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7287_ (.A0(rf_reg[343]),
    .A1(net324),
    .S(net28),
    .X(_0269_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7288_ (.A0(rf_reg[344]),
    .A1(net336),
    .S(net28),
    .X(_0270_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7289_ (.A0(rf_reg[345]),
    .A1(net333),
    .S(net27),
    .X(_0271_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7290_ (.A0(rf_reg[346]),
    .A1(net343),
    .S(net26),
    .X(_0272_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7291_ (.A0(rf_reg[347]),
    .A1(net316),
    .S(net30),
    .X(_0273_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7292_ (.A0(rf_reg[348]),
    .A1(net339),
    .S(net28),
    .X(_0274_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7293_ (.A0(rf_reg[349]),
    .A1(net335),
    .S(net26),
    .X(_0275_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7294_ (.A0(net346),
    .A1(rf_reg[34]),
    .S(net21),
    .X(_0276_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7295_ (.A0(rf_reg[350]),
    .A1(net319),
    .S(net27),
    .X(_0277_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7296_ (.A0(rf_reg[351]),
    .A1(net323),
    .S(net27),
    .X(_0278_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7297_ (.A(_2949_),
    .B(_2967_),
    .Y(_3070_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout13 (.X(net13),
    .A(net14),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7299_ (.A0(rf_reg[352]),
    .A1(net328),
    .S(net19),
    .X(_0279_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7300_ (.A0(rf_reg[353]),
    .A1(net329),
    .S(net19),
    .X(_0280_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7301_ (.A0(rf_reg[354]),
    .A1(net346),
    .S(net16),
    .X(_0281_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7302_ (.A0(rf_reg[355]),
    .A1(net331),
    .S(net20),
    .X(_0282_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7303_ (.A0(rf_reg[356]),
    .A1(net337),
    .S(net16),
    .X(_0283_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7304_ (.A0(rf_reg[357]),
    .A1(net342),
    .S(net18),
    .X(_0284_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7305_ (.A0(rf_reg[358]),
    .A1(net326),
    .S(net17),
    .X(_0285_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7306_ (.A0(rf_reg[359]),
    .A1(net340),
    .S(net18),
    .X(_0286_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7307_ (.A0(net331),
    .A1(rf_reg[35]),
    .S(net23),
    .X(_0287_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7308_ (.A0(rf_reg[360]),
    .A1(net341),
    .S(net17),
    .X(_0288_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7309_ (.A0(rf_reg[361]),
    .A1(net347),
    .S(net16),
    .X(_0289_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout12 (.X(net12),
    .A(net15),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7311_ (.A0(rf_reg[362]),
    .A1(net327),
    .S(net19),
    .X(_0290_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7312_ (.A0(rf_reg[363]),
    .A1(net317),
    .S(net19),
    .X(_0291_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7313_ (.A0(rf_reg[364]),
    .A1(net322),
    .S(net17),
    .X(_0292_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7314_ (.A0(rf_reg[365]),
    .A1(net345),
    .S(net18),
    .X(_0293_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7315_ (.A0(rf_reg[366]),
    .A1(net321),
    .S(net17),
    .X(_0294_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7316_ (.A0(rf_reg[367]),
    .A1(net332),
    .S(net19),
    .X(_0295_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7317_ (.A0(rf_reg[368]),
    .A1(net320),
    .S(net18),
    .X(_0296_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7318_ (.A0(rf_reg[369]),
    .A1(net330),
    .S(net16),
    .X(_0297_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7319_ (.A0(net337),
    .A1(rf_reg[36]),
    .S(net22),
    .X(_0298_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7320_ (.A0(rf_reg[370]),
    .A1(net318),
    .S(net19),
    .X(_0299_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7321_ (.A0(rf_reg[371]),
    .A1(net325),
    .S(net19),
    .X(_0300_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout11 (.X(net11),
    .A(net15),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7323_ (.A0(rf_reg[372]),
    .A1(net344),
    .S(net18),
    .X(_0301_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7324_ (.A0(rf_reg[373]),
    .A1(net334),
    .S(net16),
    .X(_0302_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7325_ (.A0(rf_reg[374]),
    .A1(net338),
    .S(net16),
    .X(_0303_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7326_ (.A0(rf_reg[375]),
    .A1(net324),
    .S(net18),
    .X(_0304_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7327_ (.A0(rf_reg[376]),
    .A1(net336),
    .S(net18),
    .X(_0305_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7328_ (.A0(rf_reg[377]),
    .A1(net333),
    .S(net17),
    .X(_0306_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7329_ (.A0(rf_reg[378]),
    .A1(net343),
    .S(net16),
    .X(_0307_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7330_ (.A0(rf_reg[379]),
    .A1(net316),
    .S(net20),
    .X(_0308_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7331_ (.A0(net342),
    .A1(rf_reg[37]),
    .S(net23),
    .X(_0309_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7332_ (.A0(rf_reg[380]),
    .A1(net339),
    .S(net18),
    .X(_0310_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7333_ (.A0(rf_reg[381]),
    .A1(net335),
    .S(net16),
    .X(_0311_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7334_ (.A0(rf_reg[382]),
    .A1(net319),
    .S(net17),
    .X(_0312_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7335_ (.A0(rf_reg[383]),
    .A1(net323),
    .S(net17),
    .X(_0313_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7336_ (.A(_3019_),
    .B(_3049_),
    .Y(_3074_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout10 (.X(net10),
    .A(_3078_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7338_ (.A0(rf_reg[384]),
    .A1(net328),
    .S(net14),
    .X(_0314_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7339_ (.A0(rf_reg[385]),
    .A1(net329),
    .S(net14),
    .X(_0315_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7340_ (.A0(rf_reg[386]),
    .A1(net346),
    .S(net11),
    .X(_0316_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7341_ (.A0(rf_reg[387]),
    .A1(net331),
    .S(net13),
    .X(_0317_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7342_ (.A0(rf_reg[388]),
    .A1(net337),
    .S(net11),
    .X(_0318_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7343_ (.A0(rf_reg[389]),
    .A1(net342),
    .S(net13),
    .X(_0319_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7344_ (.A0(net326),
    .A1(rf_reg[38]),
    .S(net21),
    .X(_0320_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7345_ (.A0(rf_reg[390]),
    .A1(net326),
    .S(net12),
    .X(_0321_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7346_ (.A0(rf_reg[391]),
    .A1(net340),
    .S(net13),
    .X(_0322_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7347_ (.A0(rf_reg[392]),
    .A1(net341),
    .S(net12),
    .X(_0323_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7348_ (.A0(rf_reg[393]),
    .A1(net347),
    .S(net11),
    .X(_0324_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout9 (.X(net9),
    .A(net10),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7350_ (.A0(rf_reg[394]),
    .A1(net327),
    .S(net12),
    .X(_0325_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7351_ (.A0(rf_reg[395]),
    .A1(net317),
    .S(net14),
    .X(_0326_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7352_ (.A0(rf_reg[396]),
    .A1(net322),
    .S(net12),
    .X(_0327_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7353_ (.A0(rf_reg[397]),
    .A1(net345),
    .S(net13),
    .X(_0328_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7354_ (.A0(rf_reg[398]),
    .A1(net321),
    .S(net12),
    .X(_0329_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7355_ (.A0(rf_reg[399]),
    .A1(net332),
    .S(net14),
    .X(_0330_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7356_ (.A0(net340),
    .A1(rf_reg[39]),
    .S(net23),
    .X(_0331_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7357_ (.A0(rf_reg[400]),
    .A1(net320),
    .S(net14),
    .X(_0332_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7358_ (.A0(rf_reg[401]),
    .A1(net330),
    .S(net11),
    .X(_0333_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7359_ (.A0(rf_reg[402]),
    .A1(net318),
    .S(net14),
    .X(_0334_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7360_ (.A0(rf_reg[403]),
    .A1(net325),
    .S(net14),
    .X(_0335_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout8 (.X(net8),
    .A(net9),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7362_ (.A0(rf_reg[404]),
    .A1(net344),
    .S(net13),
    .X(_0336_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7363_ (.A0(rf_reg[405]),
    .A1(net334),
    .S(net11),
    .X(_0337_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7364_ (.A0(rf_reg[406]),
    .A1(net338),
    .S(net11),
    .X(_0338_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7365_ (.A0(rf_reg[407]),
    .A1(net324),
    .S(net13),
    .X(_0339_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7366_ (.A0(rf_reg[408]),
    .A1(net336),
    .S(net13),
    .X(_0340_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7367_ (.A0(rf_reg[409]),
    .A1(net333),
    .S(net12),
    .X(_0341_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7368_ (.A0(net341),
    .A1(rf_reg[40]),
    .S(net21),
    .X(_0342_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7369_ (.A0(rf_reg[410]),
    .A1(net343),
    .S(net11),
    .X(_0343_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7370_ (.A0(rf_reg[411]),
    .A1(net316),
    .S(net15),
    .X(_0344_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7371_ (.A0(rf_reg[412]),
    .A1(net339),
    .S(net13),
    .X(_0345_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7372_ (.A0(rf_reg[413]),
    .A1(net335),
    .S(net11),
    .X(_0346_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7373_ (.A0(rf_reg[414]),
    .A1(net319),
    .S(net12),
    .X(_0347_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7374_ (.A0(rf_reg[415]),
    .A1(net323),
    .S(net12),
    .X(_0348_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7375_ (.A(_2949_),
    .B(_3019_),
    .Y(_3078_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout7 (.X(net7),
    .A(net10),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7377_ (.A0(rf_reg[416]),
    .A1(net328),
    .S(net9),
    .X(_0349_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7378_ (.A0(rf_reg[417]),
    .A1(net329),
    .S(net9),
    .X(_0350_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7379_ (.A0(rf_reg[418]),
    .A1(net346),
    .S(net6),
    .X(_0351_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7380_ (.A0(rf_reg[419]),
    .A1(net331),
    .S(net8),
    .X(_0352_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7381_ (.A0(net347),
    .A1(rf_reg[41]),
    .S(net21),
    .X(_0353_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7382_ (.A0(rf_reg[420]),
    .A1(net337),
    .S(net6),
    .X(_0354_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7383_ (.A0(rf_reg[421]),
    .A1(net342),
    .S(net8),
    .X(_0355_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7384_ (.A0(rf_reg[422]),
    .A1(net326),
    .S(net7),
    .X(_0356_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7385_ (.A0(rf_reg[423]),
    .A1(net340),
    .S(net8),
    .X(_0357_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7386_ (.A0(rf_reg[424]),
    .A1(net341),
    .S(net7),
    .X(_0358_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7387_ (.A0(rf_reg[425]),
    .A1(net347),
    .S(net6),
    .X(_0359_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout6 (.X(net6),
    .A(net10),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7389_ (.A0(rf_reg[426]),
    .A1(net327),
    .S(net7),
    .X(_0360_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7390_ (.A0(rf_reg[427]),
    .A1(net317),
    .S(net9),
    .X(_0361_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7391_ (.A0(rf_reg[428]),
    .A1(net322),
    .S(net7),
    .X(_0362_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7392_ (.A0(rf_reg[429]),
    .A1(net345),
    .S(net8),
    .X(_0363_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout5 (.X(net5),
    .A(_3083_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7394_ (.A0(net327),
    .A1(rf_reg[42]),
    .S(net22),
    .X(_0364_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7395_ (.A0(rf_reg[430]),
    .A1(net321),
    .S(net7),
    .X(_0365_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7396_ (.A0(rf_reg[431]),
    .A1(net332),
    .S(net9),
    .X(_0366_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7397_ (.A0(rf_reg[432]),
    .A1(net320),
    .S(net9),
    .X(_0367_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7398_ (.A0(rf_reg[433]),
    .A1(net330),
    .S(net6),
    .X(_0368_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7399_ (.A0(rf_reg[434]),
    .A1(net318),
    .S(net9),
    .X(_0369_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7400_ (.A0(rf_reg[435]),
    .A1(net325),
    .S(net9),
    .X(_0370_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout4 (.X(net4),
    .A(net5),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7402_ (.A0(rf_reg[436]),
    .A1(net344),
    .S(net8),
    .X(_0371_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7403_ (.A0(rf_reg[437]),
    .A1(net334),
    .S(net6),
    .X(_0372_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7404_ (.A0(rf_reg[438]),
    .A1(net338),
    .S(net6),
    .X(_0373_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7405_ (.A0(rf_reg[439]),
    .A1(net324),
    .S(net10),
    .X(_0374_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7406_ (.A0(net317),
    .A1(rf_reg[43]),
    .S(net24),
    .X(_0375_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7407_ (.A0(rf_reg[440]),
    .A1(net336),
    .S(net8),
    .X(_0376_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7408_ (.A0(rf_reg[441]),
    .A1(net333),
    .S(net7),
    .X(_0377_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7409_ (.A0(rf_reg[442]),
    .A1(net343),
    .S(net6),
    .X(_0378_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7410_ (.A0(rf_reg[443]),
    .A1(net316),
    .S(net8),
    .X(_0379_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7411_ (.A0(rf_reg[444]),
    .A1(net339),
    .S(net8),
    .X(_0380_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7412_ (.A0(rf_reg[445]),
    .A1(net335),
    .S(net6),
    .X(_0381_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7413_ (.A0(rf_reg[446]),
    .A1(net319),
    .S(net7),
    .X(_0382_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7414_ (.A0(rf_reg[447]),
    .A1(net323),
    .S(net7),
    .X(_0383_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _7415_ (.A(_3037_),
    .B(_3049_),
    .Y(_3083_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout3 (.X(net3),
    .A(net4),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7417_ (.A0(rf_reg[448]),
    .A1(net328),
    .S(net4),
    .X(_0384_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7418_ (.A0(rf_reg[449]),
    .A1(net329),
    .S(net4),
    .X(_0385_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7419_ (.A0(net322),
    .A1(rf_reg[44]),
    .S(net22),
    .X(_0386_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7420_ (.A0(rf_reg[450]),
    .A1(net346),
    .S(net1),
    .X(_0387_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7421_ (.A0(rf_reg[451]),
    .A1(net331),
    .S(net3),
    .X(_0388_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7422_ (.A0(rf_reg[452]),
    .A1(net337),
    .S(net1),
    .X(_0389_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7423_ (.A0(rf_reg[453]),
    .A1(net342),
    .S(net3),
    .X(_0390_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7424_ (.A0(rf_reg[454]),
    .A1(net326),
    .S(net2),
    .X(_0391_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7425_ (.A0(rf_reg[455]),
    .A1(net340),
    .S(net3),
    .X(_0392_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7426_ (.A0(rf_reg[456]),
    .A1(net341),
    .S(net1),
    .X(_0393_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7427_ (.A0(rf_reg[457]),
    .A1(net347),
    .S(net1),
    .X(_0394_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout2 (.X(net2),
    .A(net5),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7429_ (.A0(rf_reg[458]),
    .A1(net327),
    .S(net2),
    .X(_0395_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7430_ (.A0(rf_reg[459]),
    .A1(net317),
    .S(net4),
    .X(_0396_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7431_ (.A0(net345),
    .A1(rf_reg[45]),
    .S(net23),
    .X(_0397_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7432_ (.A0(rf_reg[460]),
    .A1(net322),
    .S(net2),
    .X(_0398_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7433_ (.A0(rf_reg[461]),
    .A1(net345),
    .S(net3),
    .X(_0399_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7434_ (.A0(rf_reg[462]),
    .A1(net321),
    .S(net2),
    .X(_0400_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7435_ (.A0(rf_reg[463]),
    .A1(net332),
    .S(net4),
    .X(_0401_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7436_ (.A0(rf_reg[464]),
    .A1(net320),
    .S(net4),
    .X(_0402_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7437_ (.A0(rf_reg[465]),
    .A1(net330),
    .S(net1),
    .X(_0403_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7438_ (.A0(rf_reg[466]),
    .A1(net318),
    .S(net4),
    .X(_0404_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7439_ (.A0(rf_reg[467]),
    .A1(net325),
    .S(net4),
    .X(_0405_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout1 (.X(net1),
    .A(net2),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7441_ (.A0(rf_reg[468]),
    .A1(net344),
    .S(net3),
    .X(_0406_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7442_ (.A0(rf_reg[469]),
    .A1(net334),
    .S(net2),
    .X(_0407_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7443_ (.A0(net321),
    .A1(rf_reg[46]),
    .S(net24),
    .X(_0408_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7444_ (.A0(rf_reg[470]),
    .A1(net338),
    .S(net1),
    .X(_0409_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7445_ (.A0(rf_reg[471]),
    .A1(net324),
    .S(net5),
    .X(_0410_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7446_ (.A0(rf_reg[472]),
    .A1(net336),
    .S(net3),
    .X(_0411_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7447_ (.A0(rf_reg[473]),
    .A1(net333),
    .S(net5),
    .X(_0412_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7448_ (.A0(rf_reg[474]),
    .A1(net343),
    .S(net1),
    .X(_0413_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7449_ (.A0(rf_reg[475]),
    .A1(net316),
    .S(net3),
    .X(_0414_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _7450_ (.A0(rf_reg[476]),
    .A1(net339),
    .S(net3),
    .X(_0415_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_123_clk_i (.X(clknet_leaf_123_clk_i),
    .A(clknet_5_5__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1000]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0000_),
    .Q_N(_4188_),
    .Q(rf_reg[1000]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1001]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(_0001_),
    .Q_N(_4187_),
    .Q(rf_reg[1001]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1002]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0002_),
    .Q_N(_4186_),
    .Q(rf_reg[1002]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1003]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0003_),
    .Q_N(_4185_),
    .Q(rf_reg[1003]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1004]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0004_),
    .Q_N(_4184_),
    .Q(rf_reg[1004]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1005]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0005_),
    .Q_N(_4183_),
    .Q(rf_reg[1005]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1006]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0006_),
    .Q_N(_4182_),
    .Q(rf_reg[1006]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1007]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0007_),
    .Q_N(_4181_),
    .Q(rf_reg[1007]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1008]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0008_),
    .Q_N(_4180_),
    .Q(rf_reg[1008]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1009]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0009_),
    .Q_N(_4179_),
    .Q(rf_reg[1009]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[100]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0010_),
    .Q_N(_4178_),
    .Q(rf_reg[100]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1010]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0011_),
    .Q_N(_4177_),
    .Q(rf_reg[1010]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1011]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0012_),
    .Q_N(_4176_),
    .Q(rf_reg[1011]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1012]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0013_),
    .Q_N(_4175_),
    .Q(rf_reg[1012]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1013]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0014_),
    .Q_N(_4174_),
    .Q(rf_reg[1013]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1014]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0015_),
    .Q_N(_4173_),
    .Q(rf_reg[1014]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1015]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0016_),
    .Q_N(_4172_),
    .Q(rf_reg[1015]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1016]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0017_),
    .Q_N(_4171_),
    .Q(rf_reg[1016]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1017]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0018_),
    .Q_N(_4170_),
    .Q(rf_reg[1017]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1018]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0019_),
    .Q_N(_4169_),
    .Q(rf_reg[1018]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1019]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0020_),
    .Q_N(_4168_),
    .Q(rf_reg[1019]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[101]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0021_),
    .Q_N(_4167_),
    .Q(rf_reg[101]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1020]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0022_),
    .Q_N(_4166_),
    .Q(rf_reg[1020]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1021]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0023_),
    .Q_N(_4165_),
    .Q(rf_reg[1021]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1022]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0024_),
    .Q_N(_4164_),
    .Q(rf_reg[1022]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[1023]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0025_),
    .Q_N(_4163_),
    .Q(rf_reg[1023]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[102]_reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(rst_ni),
    .D(_0026_),
    .Q_N(_4162_),
    .Q(rf_reg[102]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[103]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0027_),
    .Q_N(_4161_),
    .Q(rf_reg[103]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[104]_reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(rst_ni),
    .D(_0028_),
    .Q_N(_4160_),
    .Q(rf_reg[104]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[105]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0029_),
    .Q_N(_4159_),
    .Q(rf_reg[105]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[106]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0030_),
    .Q_N(_4158_),
    .Q(rf_reg[106]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[107]_reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(rst_ni),
    .D(_0031_),
    .Q_N(_4157_),
    .Q(rf_reg[107]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[108]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0032_),
    .Q_N(_4156_),
    .Q(rf_reg[108]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[109]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0033_),
    .Q_N(_4155_),
    .Q(rf_reg[109]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[110]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0034_),
    .Q_N(_4154_),
    .Q(rf_reg[110]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[111]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0035_),
    .Q_N(_4153_),
    .Q(rf_reg[111]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[112]_reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(rst_ni),
    .D(_0036_),
    .Q_N(_4152_),
    .Q(rf_reg[112]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[113]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0037_),
    .Q_N(_4151_),
    .Q(rf_reg[113]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[114]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0038_),
    .Q_N(_4150_),
    .Q(rf_reg[114]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[115]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0039_),
    .Q_N(_4149_),
    .Q(rf_reg[115]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[116]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0040_),
    .Q_N(_4148_),
    .Q(rf_reg[116]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[117]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0041_),
    .Q_N(_4147_),
    .Q(rf_reg[117]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[118]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0042_),
    .Q_N(_4146_),
    .Q(rf_reg[118]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[119]_reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(rst_ni),
    .D(_0043_),
    .Q_N(_4145_),
    .Q(rf_reg[119]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[120]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0044_),
    .Q_N(_4144_),
    .Q(rf_reg[120]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[121]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0045_),
    .Q_N(_4143_),
    .Q(rf_reg[121]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[122]_reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(rst_ni),
    .D(_0046_),
    .Q_N(_4142_),
    .Q(rf_reg[122]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[123]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0047_),
    .Q_N(_4141_),
    .Q(rf_reg[123]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[124]_reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(rst_ni),
    .D(_0048_),
    .Q_N(_4140_),
    .Q(rf_reg[124]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[125]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0049_),
    .Q_N(_4139_),
    .Q(rf_reg[125]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[126]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0050_),
    .Q_N(_4138_),
    .Q(rf_reg[126]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[127]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0051_),
    .Q_N(_4137_),
    .Q(rf_reg[127]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[128]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0052_),
    .Q_N(_4136_),
    .Q(rf_reg[128]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[129]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0053_),
    .Q_N(_4135_),
    .Q(rf_reg[129]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[130]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0054_),
    .Q_N(_4134_),
    .Q(rf_reg[130]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[131]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0055_),
    .Q_N(_4133_),
    .Q(rf_reg[131]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[132]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0056_),
    .Q_N(_4132_),
    .Q(rf_reg[132]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[133]_reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(rst_ni),
    .D(_0057_),
    .Q_N(_4131_),
    .Q(rf_reg[133]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[134]_reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(rst_ni),
    .D(_0058_),
    .Q_N(_4130_),
    .Q(rf_reg[134]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[135]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0059_),
    .Q_N(_4129_),
    .Q(rf_reg[135]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[136]_reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(rst_ni),
    .D(_0060_),
    .Q_N(_4128_),
    .Q(rf_reg[136]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[137]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0061_),
    .Q_N(_4127_),
    .Q(rf_reg[137]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[138]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0062_),
    .Q_N(_4126_),
    .Q(rf_reg[138]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[139]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0063_),
    .Q_N(_4125_),
    .Q(rf_reg[139]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[140]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0064_),
    .Q_N(_4124_),
    .Q(rf_reg[140]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[141]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0065_),
    .Q_N(_4123_),
    .Q(rf_reg[141]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[142]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0066_),
    .Q_N(_4122_),
    .Q(rf_reg[142]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[143]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0067_),
    .Q_N(_4121_),
    .Q(rf_reg[143]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[144]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0068_),
    .Q_N(_4120_),
    .Q(rf_reg[144]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[145]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0069_),
    .Q_N(_4119_),
    .Q(rf_reg[145]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[146]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0070_),
    .Q_N(_4118_),
    .Q(rf_reg[146]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[147]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0071_),
    .Q_N(_4117_),
    .Q(rf_reg[147]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[148]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0072_),
    .Q_N(_4116_),
    .Q(rf_reg[148]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[149]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0073_),
    .Q_N(_4115_),
    .Q(rf_reg[149]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[150]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0074_),
    .Q_N(_4114_),
    .Q(rf_reg[150]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[151]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0075_),
    .Q_N(_4113_),
    .Q(rf_reg[151]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[152]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0076_),
    .Q_N(_4112_),
    .Q(rf_reg[152]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[153]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0077_),
    .Q_N(_4111_),
    .Q(rf_reg[153]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[154]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0078_),
    .Q_N(_4110_),
    .Q(rf_reg[154]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[155]_reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(rst_ni),
    .D(_0079_),
    .Q_N(_4109_),
    .Q(rf_reg[155]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[156]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0080_),
    .Q_N(_4108_),
    .Q(rf_reg[156]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[157]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0081_),
    .Q_N(_4107_),
    .Q(rf_reg[157]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[158]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0082_),
    .Q_N(_4106_),
    .Q(rf_reg[158]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[159]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0083_),
    .Q_N(_4105_),
    .Q(rf_reg[159]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[160]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0084_),
    .Q_N(_4104_),
    .Q(rf_reg[160]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[161]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0085_),
    .Q_N(_4103_),
    .Q(rf_reg[161]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[162]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0086_),
    .Q_N(_4102_),
    .Q(rf_reg[162]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[163]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0087_),
    .Q_N(_4101_),
    .Q(rf_reg[163]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[164]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0088_),
    .Q_N(_4100_),
    .Q(rf_reg[164]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[165]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0089_),
    .Q_N(_4099_),
    .Q(rf_reg[165]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[166]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0090_),
    .Q_N(_4098_),
    .Q(rf_reg[166]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[167]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0091_),
    .Q_N(_4097_),
    .Q(rf_reg[167]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[168]_reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(rst_ni),
    .D(_0092_),
    .Q_N(_4096_),
    .Q(rf_reg[168]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[169]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0093_),
    .Q_N(_4095_),
    .Q(rf_reg[169]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[170]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0094_),
    .Q_N(_4094_),
    .Q(rf_reg[170]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[171]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0095_),
    .Q_N(_4093_),
    .Q(rf_reg[171]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[172]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0096_),
    .Q_N(_4092_),
    .Q(rf_reg[172]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[173]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0097_),
    .Q_N(_4091_),
    .Q(rf_reg[173]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[174]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0098_),
    .Q_N(_4090_),
    .Q(rf_reg[174]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[175]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0099_),
    .Q_N(_4089_),
    .Q(rf_reg[175]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[176]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0100_),
    .Q_N(_4088_),
    .Q(rf_reg[176]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[177]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0101_),
    .Q_N(_4087_),
    .Q(rf_reg[177]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[178]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0102_),
    .Q_N(_4086_),
    .Q(rf_reg[178]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[179]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0103_),
    .Q_N(_4085_),
    .Q(rf_reg[179]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[180]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0104_),
    .Q_N(_4084_),
    .Q(rf_reg[180]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[181]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0105_),
    .Q_N(_4083_),
    .Q(rf_reg[181]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[182]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0106_),
    .Q_N(_4082_),
    .Q(rf_reg[182]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[183]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0107_),
    .Q_N(_4081_),
    .Q(rf_reg[183]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[184]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0108_),
    .Q_N(_4080_),
    .Q(rf_reg[184]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[185]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0109_),
    .Q_N(_4079_),
    .Q(rf_reg[185]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[186]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0110_),
    .Q_N(_4078_),
    .Q(rf_reg[186]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[187]_reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(rst_ni),
    .D(_0111_),
    .Q_N(_4077_),
    .Q(rf_reg[187]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[188]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0112_),
    .Q_N(_4076_),
    .Q(rf_reg[188]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[189]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0113_),
    .Q_N(_4075_),
    .Q(rf_reg[189]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[190]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0114_),
    .Q_N(_4074_),
    .Q(rf_reg[190]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[191]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0115_),
    .Q_N(_4073_),
    .Q(rf_reg[191]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[192]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0116_),
    .Q_N(_4072_),
    .Q(rf_reg[192]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[193]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0117_),
    .Q_N(_4071_),
    .Q(rf_reg[193]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[194]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0118_),
    .Q_N(_4070_),
    .Q(rf_reg[194]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[195]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0119_),
    .Q_N(_4069_),
    .Q(rf_reg[195]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[196]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0120_),
    .Q_N(_4068_),
    .Q(rf_reg[196]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[197]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0121_),
    .Q_N(_4067_),
    .Q(rf_reg[197]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[198]_reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(rst_ni),
    .D(_0122_),
    .Q_N(_4066_),
    .Q(rf_reg[198]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[199]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0123_),
    .Q_N(_4065_),
    .Q(rf_reg[199]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[200]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0124_),
    .Q_N(_4064_),
    .Q(rf_reg[200]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[201]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0125_),
    .Q_N(_4063_),
    .Q(rf_reg[201]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[202]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0126_),
    .Q_N(_4062_),
    .Q(rf_reg[202]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[203]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0127_),
    .Q_N(_4061_),
    .Q(rf_reg[203]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[204]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0128_),
    .Q_N(_4060_),
    .Q(rf_reg[204]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[205]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0129_),
    .Q_N(_4059_),
    .Q(rf_reg[205]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[206]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0130_),
    .Q_N(_4058_),
    .Q(rf_reg[206]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[207]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0131_),
    .Q_N(_4057_),
    .Q(rf_reg[207]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[208]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0132_),
    .Q_N(_4056_),
    .Q(rf_reg[208]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[209]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0133_),
    .Q_N(_4055_),
    .Q(rf_reg[209]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[210]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0134_),
    .Q_N(_4054_),
    .Q(rf_reg[210]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[211]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0135_),
    .Q_N(_4053_),
    .Q(rf_reg[211]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[212]_reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(rst_ni),
    .D(_0136_),
    .Q_N(_4052_),
    .Q(rf_reg[212]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[213]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0137_),
    .Q_N(_4051_),
    .Q(rf_reg[213]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[214]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0138_),
    .Q_N(_4050_),
    .Q(rf_reg[214]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[215]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0139_),
    .Q_N(_4049_),
    .Q(rf_reg[215]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[216]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0140_),
    .Q_N(_4048_),
    .Q(rf_reg[216]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[217]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0141_),
    .Q_N(_4047_),
    .Q(rf_reg[217]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[218]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0142_),
    .Q_N(_4046_),
    .Q(rf_reg[218]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[219]_reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(rst_ni),
    .D(_0143_),
    .Q_N(_4045_),
    .Q(rf_reg[219]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[220]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0144_),
    .Q_N(_4044_),
    .Q(rf_reg[220]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[221]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0145_),
    .Q_N(_4043_),
    .Q(rf_reg[221]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[222]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0146_),
    .Q_N(_4042_),
    .Q(rf_reg[222]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[223]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0147_),
    .Q_N(_4041_),
    .Q(rf_reg[223]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[224]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0148_),
    .Q_N(_4040_),
    .Q(rf_reg[224]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[225]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0149_),
    .Q_N(_4039_),
    .Q(rf_reg[225]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[226]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0150_),
    .Q_N(_4038_),
    .Q(rf_reg[226]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[227]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0151_),
    .Q_N(_4037_),
    .Q(rf_reg[227]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[228]_reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(rst_ni),
    .D(_0152_),
    .Q_N(_4036_),
    .Q(rf_reg[228]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[229]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0153_),
    .Q_N(_4035_),
    .Q(rf_reg[229]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[230]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0154_),
    .Q_N(_4034_),
    .Q(rf_reg[230]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[231]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0155_),
    .Q_N(_4033_),
    .Q(rf_reg[231]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[232]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0156_),
    .Q_N(_4032_),
    .Q(rf_reg[232]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[233]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0157_),
    .Q_N(_4031_),
    .Q(rf_reg[233]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[234]_reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(rst_ni),
    .D(_0158_),
    .Q_N(_4030_),
    .Q(rf_reg[234]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[235]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0159_),
    .Q_N(_4029_),
    .Q(rf_reg[235]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[236]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0160_),
    .Q_N(_4028_),
    .Q(rf_reg[236]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[237]_reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(rst_ni),
    .D(_0161_),
    .Q_N(_4027_),
    .Q(rf_reg[237]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[238]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0162_),
    .Q_N(_4026_),
    .Q(rf_reg[238]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[239]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0163_),
    .Q_N(_4025_),
    .Q(rf_reg[239]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[240]_reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(rst_ni),
    .D(_0164_),
    .Q_N(_4024_),
    .Q(rf_reg[240]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[241]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0165_),
    .Q_N(_4023_),
    .Q(rf_reg[241]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[242]_reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(rst_ni),
    .D(_0166_),
    .Q_N(_4022_),
    .Q(rf_reg[242]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[243]_reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(rst_ni),
    .D(_0167_),
    .Q_N(_4021_),
    .Q(rf_reg[243]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[244]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0168_),
    .Q_N(_4020_),
    .Q(rf_reg[244]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[245]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0169_),
    .Q_N(_4019_),
    .Q(rf_reg[245]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[246]_reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(rst_ni),
    .D(_0170_),
    .Q_N(_4018_),
    .Q(rf_reg[246]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[247]_reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(rst_ni),
    .D(_0171_),
    .Q_N(_4017_),
    .Q(rf_reg[247]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[248]_reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(rst_ni),
    .D(_0172_),
    .Q_N(_4016_),
    .Q(rf_reg[248]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[249]_reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(rst_ni),
    .D(_0173_),
    .Q_N(_4015_),
    .Q(rf_reg[249]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[250]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0174_),
    .Q_N(_4014_),
    .Q(rf_reg[250]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[251]_reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(rst_ni),
    .D(_0175_),
    .Q_N(_4013_),
    .Q(rf_reg[251]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[252]_reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(rst_ni),
    .D(_0176_),
    .Q_N(_4012_),
    .Q(rf_reg[252]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[253]_reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(rst_ni),
    .D(_0177_),
    .Q_N(_4011_),
    .Q(rf_reg[253]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[254]_reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(rst_ni),
    .D(_0178_),
    .Q_N(_4010_),
    .Q(rf_reg[254]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[255]_reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(rst_ni),
    .D(_0179_),
    .Q_N(_4009_),
    .Q(rf_reg[255]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[256]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0180_),
    .Q_N(_4008_),
    .Q(rf_reg[256]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[257]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0181_),
    .Q_N(_4007_),
    .Q(rf_reg[257]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[258]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0182_),
    .Q_N(_4006_),
    .Q(rf_reg[258]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[259]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0183_),
    .Q_N(_4005_),
    .Q(rf_reg[259]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[260]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0184_),
    .Q_N(_4004_),
    .Q(rf_reg[260]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[261]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0185_),
    .Q_N(_4003_),
    .Q(rf_reg[261]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[262]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0186_),
    .Q_N(_4002_),
    .Q(rf_reg[262]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[263]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0187_),
    .Q_N(_4001_),
    .Q(rf_reg[263]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[264]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0188_),
    .Q_N(_4000_),
    .Q(rf_reg[264]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[265]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0189_),
    .Q_N(_3999_),
    .Q(rf_reg[265]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[266]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0190_),
    .Q_N(_3998_),
    .Q(rf_reg[266]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[267]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0191_),
    .Q_N(_3997_),
    .Q(rf_reg[267]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[268]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0192_),
    .Q_N(_3996_),
    .Q(rf_reg[268]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[269]_reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(rst_ni),
    .D(_0193_),
    .Q_N(_3995_),
    .Q(rf_reg[269]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[270]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0194_),
    .Q_N(_3994_),
    .Q(rf_reg[270]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[271]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0195_),
    .Q_N(_3993_),
    .Q(rf_reg[271]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[272]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0196_),
    .Q_N(_3992_),
    .Q(rf_reg[272]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[273]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0197_),
    .Q_N(_3991_),
    .Q(rf_reg[273]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[274]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0198_),
    .Q_N(_3990_),
    .Q(rf_reg[274]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[275]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0199_),
    .Q_N(_3989_),
    .Q(rf_reg[275]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[276]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0200_),
    .Q_N(_3988_),
    .Q(rf_reg[276]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[277]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0201_),
    .Q_N(_3987_),
    .Q(rf_reg[277]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[278]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0202_),
    .Q_N(_3986_),
    .Q(rf_reg[278]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[279]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0203_),
    .Q_N(_3985_),
    .Q(rf_reg[279]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[280]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0204_),
    .Q_N(_3984_),
    .Q(rf_reg[280]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[281]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0205_),
    .Q_N(_3983_),
    .Q(rf_reg[281]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[282]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0206_),
    .Q_N(_3982_),
    .Q(rf_reg[282]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[283]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0207_),
    .Q_N(_3981_),
    .Q(rf_reg[283]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[284]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0208_),
    .Q_N(_3980_),
    .Q(rf_reg[284]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[285]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0209_),
    .Q_N(_3979_),
    .Q(rf_reg[285]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[286]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0210_),
    .Q_N(_3978_),
    .Q(rf_reg[286]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[287]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0211_),
    .Q_N(_3977_),
    .Q(rf_reg[287]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[288]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0212_),
    .Q_N(_3976_),
    .Q(rf_reg[288]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[289]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0213_),
    .Q_N(_3975_),
    .Q(rf_reg[289]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[290]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0214_),
    .Q_N(_3974_),
    .Q(rf_reg[290]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[291]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0215_),
    .Q_N(_3973_),
    .Q(rf_reg[291]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[292]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0216_),
    .Q_N(_3972_),
    .Q(rf_reg[292]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[293]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0217_),
    .Q_N(_3971_),
    .Q(rf_reg[293]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[294]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0218_),
    .Q_N(_3970_),
    .Q(rf_reg[294]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[295]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0219_),
    .Q_N(_3969_),
    .Q(rf_reg[295]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[296]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0220_),
    .Q_N(_3968_),
    .Q(rf_reg[296]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[297]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0221_),
    .Q_N(_3967_),
    .Q(rf_reg[297]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[298]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0222_),
    .Q_N(_3966_),
    .Q(rf_reg[298]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[299]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0223_),
    .Q_N(_3965_),
    .Q(rf_reg[299]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[300]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0224_),
    .Q_N(_3964_),
    .Q(rf_reg[300]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[301]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0225_),
    .Q_N(_3963_),
    .Q(rf_reg[301]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[302]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0226_),
    .Q_N(_3962_),
    .Q(rf_reg[302]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[303]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0227_),
    .Q_N(_3961_),
    .Q(rf_reg[303]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[304]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0228_),
    .Q_N(_3960_),
    .Q(rf_reg[304]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[305]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0229_),
    .Q_N(_3959_),
    .Q(rf_reg[305]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[306]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0230_),
    .Q_N(_3958_),
    .Q(rf_reg[306]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[307]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0231_),
    .Q_N(_3957_),
    .Q(rf_reg[307]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[308]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0232_),
    .Q_N(_3956_),
    .Q(rf_reg[308]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[309]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0233_),
    .Q_N(_3955_),
    .Q(rf_reg[309]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[310]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0234_),
    .Q_N(_3954_),
    .Q(rf_reg[310]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[311]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0235_),
    .Q_N(_3953_),
    .Q(rf_reg[311]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[312]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0236_),
    .Q_N(_3952_),
    .Q(rf_reg[312]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[313]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0237_),
    .Q_N(_3951_),
    .Q(rf_reg[313]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[314]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0238_),
    .Q_N(_3950_),
    .Q(rf_reg[314]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[315]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0239_),
    .Q_N(_3949_),
    .Q(rf_reg[315]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[316]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0240_),
    .Q_N(_3948_),
    .Q(rf_reg[316]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[317]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0241_),
    .Q_N(_3947_),
    .Q(rf_reg[317]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[318]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0242_),
    .Q_N(_3946_),
    .Q(rf_reg[318]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[319]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0243_),
    .Q_N(_3945_),
    .Q(rf_reg[319]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[320]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0244_),
    .Q_N(_3944_),
    .Q(rf_reg[320]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[321]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0245_),
    .Q_N(_3943_),
    .Q(rf_reg[321]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[322]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0246_),
    .Q_N(_3942_),
    .Q(rf_reg[322]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[323]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0247_),
    .Q_N(_3941_),
    .Q(rf_reg[323]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[324]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0248_),
    .Q_N(_3940_),
    .Q(rf_reg[324]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[325]_reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(rst_ni),
    .D(_0249_),
    .Q_N(_3939_),
    .Q(rf_reg[325]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[326]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0250_),
    .Q_N(_3938_),
    .Q(rf_reg[326]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[327]_reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(rst_ni),
    .D(_0251_),
    .Q_N(_3937_),
    .Q(rf_reg[327]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[328]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0252_),
    .Q_N(_3936_),
    .Q(rf_reg[328]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[329]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0253_),
    .Q_N(_3935_),
    .Q(rf_reg[329]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[32]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0254_),
    .Q_N(_3934_),
    .Q(rf_reg[32]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[330]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0255_),
    .Q_N(_3933_),
    .Q(rf_reg[330]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[331]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0256_),
    .Q_N(_3932_),
    .Q(rf_reg[331]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[332]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0257_),
    .Q_N(_3931_),
    .Q(rf_reg[332]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[333]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0258_),
    .Q_N(_3930_),
    .Q(rf_reg[333]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[334]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0259_),
    .Q_N(_3929_),
    .Q(rf_reg[334]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[335]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0260_),
    .Q_N(_3928_),
    .Q(rf_reg[335]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[336]_reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(rst_ni),
    .D(_0261_),
    .Q_N(_3927_),
    .Q(rf_reg[336]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[337]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0262_),
    .Q_N(_3926_),
    .Q(rf_reg[337]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[338]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0263_),
    .Q_N(_3925_),
    .Q(rf_reg[338]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[339]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0264_),
    .Q_N(_3924_),
    .Q(rf_reg[339]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[33]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0265_),
    .Q_N(_3923_),
    .Q(rf_reg[33]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[340]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0266_),
    .Q_N(_3922_),
    .Q(rf_reg[340]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[341]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0267_),
    .Q_N(_3921_),
    .Q(rf_reg[341]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[342]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0268_),
    .Q_N(_3920_),
    .Q(rf_reg[342]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[343]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0269_),
    .Q_N(_3919_),
    .Q(rf_reg[343]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[344]_reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(rst_ni),
    .D(_0270_),
    .Q_N(_3918_),
    .Q(rf_reg[344]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[345]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0271_),
    .Q_N(_3917_),
    .Q(rf_reg[345]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[346]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0272_),
    .Q_N(_3916_),
    .Q(rf_reg[346]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[347]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0273_),
    .Q_N(_3915_),
    .Q(rf_reg[347]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[348]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0274_),
    .Q_N(_3914_),
    .Q(rf_reg[348]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[349]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0275_),
    .Q_N(_3913_),
    .Q(rf_reg[349]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[34]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0276_),
    .Q_N(_3912_),
    .Q(rf_reg[34]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[350]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0277_),
    .Q_N(_3911_),
    .Q(rf_reg[350]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[351]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0278_),
    .Q_N(_3910_),
    .Q(rf_reg[351]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[352]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0279_),
    .Q_N(_3909_),
    .Q(rf_reg[352]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[353]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0280_),
    .Q_N(_3908_),
    .Q(rf_reg[353]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[354]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0281_),
    .Q_N(_3907_),
    .Q(rf_reg[354]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[355]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0282_),
    .Q_N(_3906_),
    .Q(rf_reg[355]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[356]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0283_),
    .Q_N(_3905_),
    .Q(rf_reg[356]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[357]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0284_),
    .Q_N(_3904_),
    .Q(rf_reg[357]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[358]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0285_),
    .Q_N(_3903_),
    .Q(rf_reg[358]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[359]_reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(rst_ni),
    .D(_0286_),
    .Q_N(_3902_),
    .Q(rf_reg[359]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[35]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0287_),
    .Q_N(_3901_),
    .Q(rf_reg[35]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[360]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0288_),
    .Q_N(_3900_),
    .Q(rf_reg[360]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[361]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0289_),
    .Q_N(_3899_),
    .Q(rf_reg[361]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[362]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0290_),
    .Q_N(_3898_),
    .Q(rf_reg[362]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[363]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0291_),
    .Q_N(_3897_),
    .Q(rf_reg[363]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[364]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0292_),
    .Q_N(_3896_),
    .Q(rf_reg[364]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[365]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0293_),
    .Q_N(_3895_),
    .Q(rf_reg[365]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[366]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0294_),
    .Q_N(_3894_),
    .Q(rf_reg[366]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[367]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0295_),
    .Q_N(_3893_),
    .Q(rf_reg[367]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[368]_reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(rst_ni),
    .D(_0296_),
    .Q_N(_3892_),
    .Q(rf_reg[368]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[369]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0297_),
    .Q_N(_3891_),
    .Q(rf_reg[369]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[36]_reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(rst_ni),
    .D(_0298_),
    .Q_N(_3890_),
    .Q(rf_reg[36]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[370]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0299_),
    .Q_N(_3889_),
    .Q(rf_reg[370]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[371]_reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(rst_ni),
    .D(_0300_),
    .Q_N(_3888_),
    .Q(rf_reg[371]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[372]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0301_),
    .Q_N(_3887_),
    .Q(rf_reg[372]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[373]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0302_),
    .Q_N(_3886_),
    .Q(rf_reg[373]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[374]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0303_),
    .Q_N(_3885_),
    .Q(rf_reg[374]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[375]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0304_),
    .Q_N(_3884_),
    .Q(rf_reg[375]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[376]_reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(rst_ni),
    .D(_0305_),
    .Q_N(_3883_),
    .Q(rf_reg[376]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[377]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0306_),
    .Q_N(_3882_),
    .Q(rf_reg[377]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[378]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0307_),
    .Q_N(_3881_),
    .Q(rf_reg[378]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[379]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0308_),
    .Q_N(_3880_),
    .Q(rf_reg[379]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[37]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0309_),
    .Q_N(_3879_),
    .Q(rf_reg[37]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[380]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(rst_ni),
    .D(_0310_),
    .Q_N(_3878_),
    .Q(rf_reg[380]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[381]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0311_),
    .Q_N(_3877_),
    .Q(rf_reg[381]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[382]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0312_),
    .Q_N(_3876_),
    .Q(rf_reg[382]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[383]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0313_),
    .Q_N(_3875_),
    .Q(rf_reg[383]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[384]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0314_),
    .Q_N(_3874_),
    .Q(rf_reg[384]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[385]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0315_),
    .Q_N(_3873_),
    .Q(rf_reg[385]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[386]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0316_),
    .Q_N(_3872_),
    .Q(rf_reg[386]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[387]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0317_),
    .Q_N(_3871_),
    .Q(rf_reg[387]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[388]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0318_),
    .Q_N(_3870_),
    .Q(rf_reg[388]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[389]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0319_),
    .Q_N(_3869_),
    .Q(rf_reg[389]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[38]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0320_),
    .Q_N(_3868_),
    .Q(rf_reg[38]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[390]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0321_),
    .Q_N(_3867_),
    .Q(rf_reg[390]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[391]_reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(rst_ni),
    .D(_0322_),
    .Q_N(_3866_),
    .Q(rf_reg[391]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[392]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0323_),
    .Q_N(_3865_),
    .Q(rf_reg[392]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[393]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(_0324_),
    .Q_N(_3864_),
    .Q(rf_reg[393]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[394]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0325_),
    .Q_N(_3863_),
    .Q(rf_reg[394]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[395]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0326_),
    .Q_N(_3862_),
    .Q(rf_reg[395]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[396]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0327_),
    .Q_N(_3861_),
    .Q(rf_reg[396]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[397]_reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(rst_ni),
    .D(_0328_),
    .Q_N(_3860_),
    .Q(rf_reg[397]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[398]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0329_),
    .Q_N(_3859_),
    .Q(rf_reg[398]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[399]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0330_),
    .Q_N(_3858_),
    .Q(rf_reg[399]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[39]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0331_),
    .Q_N(_3857_),
    .Q(rf_reg[39]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[400]_reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(rst_ni),
    .D(_0332_),
    .Q_N(_3856_),
    .Q(rf_reg[400]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[401]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0333_),
    .Q_N(_3855_),
    .Q(rf_reg[401]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[402]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0334_),
    .Q_N(_3854_),
    .Q(rf_reg[402]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[403]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0335_),
    .Q_N(_3853_),
    .Q(rf_reg[403]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[404]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0336_),
    .Q_N(_3852_),
    .Q(rf_reg[404]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[405]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0337_),
    .Q_N(_3851_),
    .Q(rf_reg[405]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[406]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0338_),
    .Q_N(_3850_),
    .Q(rf_reg[406]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[407]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0339_),
    .Q_N(_3849_),
    .Q(rf_reg[407]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[408]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0340_),
    .Q_N(_3848_),
    .Q(rf_reg[408]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[409]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0341_),
    .Q_N(_3847_),
    .Q(rf_reg[409]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[40]_reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(rst_ni),
    .D(_0342_),
    .Q_N(_3846_),
    .Q(rf_reg[40]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[410]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0343_),
    .Q_N(_3845_),
    .Q(rf_reg[410]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[411]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0344_),
    .Q_N(_3844_),
    .Q(rf_reg[411]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[412]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0345_),
    .Q_N(_3843_),
    .Q(rf_reg[412]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[413]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0346_),
    .Q_N(_3842_),
    .Q(rf_reg[413]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[414]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0347_),
    .Q_N(_3841_),
    .Q(rf_reg[414]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[415]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0348_),
    .Q_N(_3840_),
    .Q(rf_reg[415]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[416]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0349_),
    .Q_N(_3839_),
    .Q(rf_reg[416]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[417]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0350_),
    .Q_N(_3838_),
    .Q(rf_reg[417]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[418]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0351_),
    .Q_N(_3837_),
    .Q(rf_reg[418]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[419]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0352_),
    .Q_N(_3836_),
    .Q(rf_reg[419]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[41]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0353_),
    .Q_N(_3835_),
    .Q(rf_reg[41]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[420]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0354_),
    .Q_N(_3834_),
    .Q(rf_reg[420]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[421]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0355_),
    .Q_N(_3833_),
    .Q(rf_reg[421]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[422]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0356_),
    .Q_N(_3832_),
    .Q(rf_reg[422]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[423]_reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(rst_ni),
    .D(_0357_),
    .Q_N(_3831_),
    .Q(rf_reg[423]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[424]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0358_),
    .Q_N(_3830_),
    .Q(rf_reg[424]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[425]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0359_),
    .Q_N(_3829_),
    .Q(rf_reg[425]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[426]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0360_),
    .Q_N(_3828_),
    .Q(rf_reg[426]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[427]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0361_),
    .Q_N(_3827_),
    .Q(rf_reg[427]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[428]_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(rst_ni),
    .D(_0362_),
    .Q_N(_3826_),
    .Q(rf_reg[428]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[429]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0363_),
    .Q_N(_3825_),
    .Q(rf_reg[429]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[42]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0364_),
    .Q_N(_3824_),
    .Q(rf_reg[42]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[430]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0365_),
    .Q_N(_3823_),
    .Q(rf_reg[430]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[431]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0366_),
    .Q_N(_3822_),
    .Q(rf_reg[431]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[432]_reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(rst_ni),
    .D(_0367_),
    .Q_N(_3821_),
    .Q(rf_reg[432]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[433]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0368_),
    .Q_N(_3820_),
    .Q(rf_reg[433]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[434]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0369_),
    .Q_N(_3819_),
    .Q(rf_reg[434]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[435]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0370_),
    .Q_N(_3818_),
    .Q(rf_reg[435]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[436]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0371_),
    .Q_N(_3817_),
    .Q(rf_reg[436]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[437]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0372_),
    .Q_N(_3816_),
    .Q(rf_reg[437]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[438]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0373_),
    .Q_N(_3815_),
    .Q(rf_reg[438]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[439]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0374_),
    .Q_N(_3814_),
    .Q(rf_reg[439]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[43]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0375_),
    .Q_N(_3813_),
    .Q(rf_reg[43]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[440]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0376_),
    .Q_N(_3812_),
    .Q(rf_reg[440]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[441]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0377_),
    .Q_N(_3811_),
    .Q(rf_reg[441]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[442]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0378_),
    .Q_N(_3810_),
    .Q(rf_reg[442]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[443]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0379_),
    .Q_N(_3809_),
    .Q(rf_reg[443]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[444]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0380_),
    .Q_N(_3808_),
    .Q(rf_reg[444]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[445]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0381_),
    .Q_N(_3807_),
    .Q(rf_reg[445]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[446]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0382_),
    .Q_N(_3806_),
    .Q(rf_reg[446]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[447]_reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(rst_ni),
    .D(_0383_),
    .Q_N(_3805_),
    .Q(rf_reg[447]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[448]_reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(rst_ni),
    .D(_0384_),
    .Q_N(_3804_),
    .Q(rf_reg[448]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[449]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0385_),
    .Q_N(_3803_),
    .Q(rf_reg[449]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[44]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0386_),
    .Q_N(_3802_),
    .Q(rf_reg[44]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[450]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0387_),
    .Q_N(_3801_),
    .Q(rf_reg[450]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[451]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0388_),
    .Q_N(_3800_),
    .Q(rf_reg[451]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[452]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0389_),
    .Q_N(_3799_),
    .Q(rf_reg[452]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[453]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0390_),
    .Q_N(_3798_),
    .Q(rf_reg[453]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[454]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0391_),
    .Q_N(_3797_),
    .Q(rf_reg[454]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[455]_reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(rst_ni),
    .D(_0392_),
    .Q_N(_3796_),
    .Q(rf_reg[455]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[456]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0393_),
    .Q_N(_3795_),
    .Q(rf_reg[456]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[457]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0394_),
    .Q_N(_3794_),
    .Q(rf_reg[457]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[458]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0395_),
    .Q_N(_3793_),
    .Q(rf_reg[458]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[459]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0396_),
    .Q_N(_3792_),
    .Q(rf_reg[459]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[45]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0397_),
    .Q_N(_3791_),
    .Q(rf_reg[45]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[460]_reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(rst_ni),
    .D(_0398_),
    .Q_N(_3790_),
    .Q(rf_reg[460]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[461]_reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(rst_ni),
    .D(_0399_),
    .Q_N(_3789_),
    .Q(rf_reg[461]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[462]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0400_),
    .Q_N(_3788_),
    .Q(rf_reg[462]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[463]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0401_),
    .Q_N(_3787_),
    .Q(rf_reg[463]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[464]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0402_),
    .Q_N(_3786_),
    .Q(rf_reg[464]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[465]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0403_),
    .Q_N(_3785_),
    .Q(rf_reg[465]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[466]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0404_),
    .Q_N(_3784_),
    .Q(rf_reg[466]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[467]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0405_),
    .Q_N(_3783_),
    .Q(rf_reg[467]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[468]_reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(rst_ni),
    .D(_0406_),
    .Q_N(_3782_),
    .Q(rf_reg[468]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[469]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0407_),
    .Q_N(_3781_),
    .Q(rf_reg[469]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[46]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0408_),
    .Q_N(_3780_),
    .Q(rf_reg[46]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[470]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0409_),
    .Q_N(_3779_),
    .Q(rf_reg[470]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[471]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0410_),
    .Q_N(_3778_),
    .Q(rf_reg[471]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[472]_reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(rst_ni),
    .D(_0411_),
    .Q_N(_3777_),
    .Q(rf_reg[472]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[473]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0412_),
    .Q_N(_3776_),
    .Q(rf_reg[473]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[474]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0413_),
    .Q_N(_3775_),
    .Q(rf_reg[474]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[475]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0414_),
    .Q_N(_3774_),
    .Q(rf_reg[475]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[476]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0415_),
    .Q_N(_3773_),
    .Q(rf_reg[476]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[477]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0416_),
    .Q_N(_3772_),
    .Q(rf_reg[477]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[478]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0417_),
    .Q_N(_3771_),
    .Q(rf_reg[478]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[479]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0418_),
    .Q_N(_3770_),
    .Q(rf_reg[479]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[47]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0419_),
    .Q_N(_3769_),
    .Q(rf_reg[47]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[480]_reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(rst_ni),
    .D(_0420_),
    .Q_N(_3768_),
    .Q(rf_reg[480]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[481]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0421_),
    .Q_N(_3767_),
    .Q(rf_reg[481]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[482]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0422_),
    .Q_N(_3766_),
    .Q(rf_reg[482]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[483]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0423_),
    .Q_N(_3765_),
    .Q(rf_reg[483]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[484]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0424_),
    .Q_N(_3764_),
    .Q(rf_reg[484]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[485]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0425_),
    .Q_N(_3763_),
    .Q(rf_reg[485]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[486]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0426_),
    .Q_N(_3762_),
    .Q(rf_reg[486]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[487]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0427_),
    .Q_N(_3761_),
    .Q(rf_reg[487]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[488]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0428_),
    .Q_N(_3760_),
    .Q(rf_reg[488]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[489]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0429_),
    .Q_N(_3759_),
    .Q(rf_reg[489]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[48]_reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(rst_ni),
    .D(_0430_),
    .Q_N(_3758_),
    .Q(rf_reg[48]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[490]_reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(rst_ni),
    .D(_0431_),
    .Q_N(_3757_),
    .Q(rf_reg[490]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[491]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0432_),
    .Q_N(_3756_),
    .Q(rf_reg[491]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[492]_reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(rst_ni),
    .D(_0433_),
    .Q_N(_3755_),
    .Q(rf_reg[492]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[493]_reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(rst_ni),
    .D(_0434_),
    .Q_N(_3754_),
    .Q(rf_reg[493]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[494]_reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(rst_ni),
    .D(_0435_),
    .Q_N(_3753_),
    .Q(rf_reg[494]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[495]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0436_),
    .Q_N(_3752_),
    .Q(rf_reg[495]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[496]_reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(rst_ni),
    .D(_0437_),
    .Q_N(_3751_),
    .Q(rf_reg[496]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[497]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0438_),
    .Q_N(_3750_),
    .Q(rf_reg[497]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[498]_reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(rst_ni),
    .D(_0439_),
    .Q_N(_3749_),
    .Q(rf_reg[498]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[499]_reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(rst_ni),
    .D(_0440_),
    .Q_N(_3748_),
    .Q(rf_reg[499]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[49]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0441_),
    .Q_N(_3747_),
    .Q(rf_reg[49]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[500]_reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(rst_ni),
    .D(_0442_),
    .Q_N(_3746_),
    .Q(rf_reg[500]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[501]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0443_),
    .Q_N(_3745_),
    .Q(rf_reg[501]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[502]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0444_),
    .Q_N(_3744_),
    .Q(rf_reg[502]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[503]_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(rst_ni),
    .D(_0445_),
    .Q_N(_3743_),
    .Q(rf_reg[503]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[504]_reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(rst_ni),
    .D(_0446_),
    .Q_N(_3742_),
    .Q(rf_reg[504]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[505]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0447_),
    .Q_N(_3741_),
    .Q(rf_reg[505]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[506]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0448_),
    .Q_N(_3740_),
    .Q(rf_reg[506]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[507]_reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(rst_ni),
    .D(_0449_),
    .Q_N(_3739_),
    .Q(rf_reg[507]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[508]_reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(rst_ni),
    .D(_0450_),
    .Q_N(_3738_),
    .Q(rf_reg[508]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[509]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0451_),
    .Q_N(_3737_),
    .Q(rf_reg[509]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[50]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0452_),
    .Q_N(_3736_),
    .Q(rf_reg[50]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[510]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0453_),
    .Q_N(_3735_),
    .Q(rf_reg[510]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[511]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0454_),
    .Q_N(_3734_),
    .Q(rf_reg[511]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[512]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0455_),
    .Q_N(_3733_),
    .Q(rf_reg[512]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[513]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0456_),
    .Q_N(_3732_),
    .Q(rf_reg[513]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[514]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0457_),
    .Q_N(_3731_),
    .Q(rf_reg[514]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[515]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0458_),
    .Q_N(_3730_),
    .Q(rf_reg[515]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[516]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0459_),
    .Q_N(_3729_),
    .Q(rf_reg[516]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[517]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0460_),
    .Q_N(_3728_),
    .Q(rf_reg[517]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[518]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0461_),
    .Q_N(_3727_),
    .Q(rf_reg[518]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[519]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0462_),
    .Q_N(_3726_),
    .Q(rf_reg[519]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[51]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0463_),
    .Q_N(_3725_),
    .Q(rf_reg[51]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[520]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0464_),
    .Q_N(_3724_),
    .Q(rf_reg[520]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[521]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0465_),
    .Q_N(_3723_),
    .Q(rf_reg[521]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[522]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0466_),
    .Q_N(_3722_),
    .Q(rf_reg[522]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[523]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0467_),
    .Q_N(_3721_),
    .Q(rf_reg[523]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[524]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0468_),
    .Q_N(_3720_),
    .Q(rf_reg[524]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[525]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0469_),
    .Q_N(_3719_),
    .Q(rf_reg[525]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[526]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0470_),
    .Q_N(_3718_),
    .Q(rf_reg[526]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[527]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0471_),
    .Q_N(_3717_),
    .Q(rf_reg[527]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[528]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0472_),
    .Q_N(_3716_),
    .Q(rf_reg[528]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[529]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0473_),
    .Q_N(_3715_),
    .Q(rf_reg[529]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[52]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0474_),
    .Q_N(_3714_),
    .Q(rf_reg[52]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[530]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0475_),
    .Q_N(_3713_),
    .Q(rf_reg[530]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[531]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0476_),
    .Q_N(_3712_),
    .Q(rf_reg[531]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[532]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0477_),
    .Q_N(_3711_),
    .Q(rf_reg[532]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[533]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0478_),
    .Q_N(_3710_),
    .Q(rf_reg[533]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[534]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0479_),
    .Q_N(_3709_),
    .Q(rf_reg[534]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[535]_reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(rst_ni),
    .D(_0480_),
    .Q_N(_3708_),
    .Q(rf_reg[535]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[536]_reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(rst_ni),
    .D(_0481_),
    .Q_N(_3707_),
    .Q(rf_reg[536]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[537]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0482_),
    .Q_N(_3706_),
    .Q(rf_reg[537]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[538]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(_0483_),
    .Q_N(_3705_),
    .Q(rf_reg[538]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[539]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0484_),
    .Q_N(_3704_),
    .Q(rf_reg[539]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[53]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0485_),
    .Q_N(_3703_),
    .Q(rf_reg[53]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[540]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0486_),
    .Q_N(_3702_),
    .Q(rf_reg[540]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[541]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0487_),
    .Q_N(_3701_),
    .Q(rf_reg[541]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[542]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0488_),
    .Q_N(_3700_),
    .Q(rf_reg[542]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[543]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0489_),
    .Q_N(_3699_),
    .Q(rf_reg[543]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[544]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0490_),
    .Q_N(_3698_),
    .Q(rf_reg[544]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[545]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0491_),
    .Q_N(_3697_),
    .Q(rf_reg[545]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[546]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0492_),
    .Q_N(_3696_),
    .Q(rf_reg[546]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[547]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0493_),
    .Q_N(_3695_),
    .Q(rf_reg[547]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[548]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0494_),
    .Q_N(_3694_),
    .Q(rf_reg[548]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[549]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0495_),
    .Q_N(_3693_),
    .Q(rf_reg[549]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[54]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0496_),
    .Q_N(_3692_),
    .Q(rf_reg[54]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[550]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0497_),
    .Q_N(_3691_),
    .Q(rf_reg[550]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[551]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0498_),
    .Q_N(_3690_),
    .Q(rf_reg[551]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[552]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0499_),
    .Q_N(_3689_),
    .Q(rf_reg[552]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[553]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0500_),
    .Q_N(_3688_),
    .Q(rf_reg[553]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[554]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0501_),
    .Q_N(_3687_),
    .Q(rf_reg[554]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[555]_reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(rst_ni),
    .D(_0502_),
    .Q_N(_3686_),
    .Q(rf_reg[555]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[556]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0503_),
    .Q_N(_3685_),
    .Q(rf_reg[556]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[557]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0504_),
    .Q_N(_3684_),
    .Q(rf_reg[557]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[558]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0505_),
    .Q_N(_3683_),
    .Q(rf_reg[558]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[559]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0506_),
    .Q_N(_3682_),
    .Q(rf_reg[559]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[55]_reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(rst_ni),
    .D(_0507_),
    .Q_N(_3681_),
    .Q(rf_reg[55]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[560]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0508_),
    .Q_N(_3680_),
    .Q(rf_reg[560]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[561]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0509_),
    .Q_N(_3679_),
    .Q(rf_reg[561]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[562]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0510_),
    .Q_N(_3678_),
    .Q(rf_reg[562]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[563]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0511_),
    .Q_N(_3677_),
    .Q(rf_reg[563]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[564]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0512_),
    .Q_N(_3676_),
    .Q(rf_reg[564]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[565]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0513_),
    .Q_N(_3675_),
    .Q(rf_reg[565]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[566]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0514_),
    .Q_N(_3674_),
    .Q(rf_reg[566]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[567]_reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(rst_ni),
    .D(_0515_),
    .Q_N(_3673_),
    .Q(rf_reg[567]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[568]_reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(rst_ni),
    .D(_0516_),
    .Q_N(_3672_),
    .Q(rf_reg[568]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[569]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0517_),
    .Q_N(_3671_),
    .Q(rf_reg[569]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[56]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0518_),
    .Q_N(_3670_),
    .Q(rf_reg[56]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[570]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0519_),
    .Q_N(_3669_),
    .Q(rf_reg[570]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[571]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0520_),
    .Q_N(_3668_),
    .Q(rf_reg[571]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[572]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0521_),
    .Q_N(_3667_),
    .Q(rf_reg[572]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[573]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0522_),
    .Q_N(_3666_),
    .Q(rf_reg[573]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[574]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0523_),
    .Q_N(_3665_),
    .Q(rf_reg[574]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[575]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0524_),
    .Q_N(_3664_),
    .Q(rf_reg[575]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[576]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0525_),
    .Q_N(_3663_),
    .Q(rf_reg[576]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[577]_reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(rst_ni),
    .D(_0526_),
    .Q_N(_3662_),
    .Q(rf_reg[577]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[578]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0527_),
    .Q_N(_3661_),
    .Q(rf_reg[578]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[579]_reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(rst_ni),
    .D(_0528_),
    .Q_N(_3660_),
    .Q(rf_reg[579]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[57]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0529_),
    .Q_N(_3659_),
    .Q(rf_reg[57]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[580]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0530_),
    .Q_N(_3658_),
    .Q(rf_reg[580]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[581]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0531_),
    .Q_N(_3657_),
    .Q(rf_reg[581]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[582]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0532_),
    .Q_N(_3656_),
    .Q(rf_reg[582]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[583]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0533_),
    .Q_N(_3655_),
    .Q(rf_reg[583]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[584]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0534_),
    .Q_N(_3654_),
    .Q(rf_reg[584]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[585]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0535_),
    .Q_N(_3653_),
    .Q(rf_reg[585]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[586]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0536_),
    .Q_N(_3652_),
    .Q(rf_reg[586]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[587]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0537_),
    .Q_N(_3651_),
    .Q(rf_reg[587]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[588]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0538_),
    .Q_N(_3650_),
    .Q(rf_reg[588]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[589]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0539_),
    .Q_N(_3649_),
    .Q(rf_reg[589]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[58]_reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(rst_ni),
    .D(_0540_),
    .Q_N(_3648_),
    .Q(rf_reg[58]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[590]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0541_),
    .Q_N(_3647_),
    .Q(rf_reg[590]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[591]_reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(rst_ni),
    .D(_0542_),
    .Q_N(_3646_),
    .Q(rf_reg[591]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[592]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0543_),
    .Q_N(_3645_),
    .Q(rf_reg[592]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[593]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0544_),
    .Q_N(_3644_),
    .Q(rf_reg[593]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[594]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0545_),
    .Q_N(_3643_),
    .Q(rf_reg[594]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[595]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0546_),
    .Q_N(_3642_),
    .Q(rf_reg[595]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[596]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0547_),
    .Q_N(_3641_),
    .Q(rf_reg[596]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[597]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0548_),
    .Q_N(_3640_),
    .Q(rf_reg[597]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[598]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0549_),
    .Q_N(_3639_),
    .Q(rf_reg[598]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[599]_reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(rst_ni),
    .D(_0550_),
    .Q_N(_3638_),
    .Q(rf_reg[599]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[59]_reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(rst_ni),
    .D(_0551_),
    .Q_N(_3637_),
    .Q(rf_reg[59]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[600]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0552_),
    .Q_N(_3636_),
    .Q(rf_reg[600]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[601]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0553_),
    .Q_N(_3635_),
    .Q(rf_reg[601]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[602]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(_0554_),
    .Q_N(_3634_),
    .Q(rf_reg[602]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[603]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0555_),
    .Q_N(_3633_),
    .Q(rf_reg[603]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[604]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0556_),
    .Q_N(_3632_),
    .Q(rf_reg[604]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[605]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0557_),
    .Q_N(_3631_),
    .Q(rf_reg[605]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[606]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0558_),
    .Q_N(_3630_),
    .Q(rf_reg[606]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[607]_reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(rst_ni),
    .D(_0559_),
    .Q_N(_3629_),
    .Q(rf_reg[607]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[608]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0560_),
    .Q_N(_3628_),
    .Q(rf_reg[608]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[609]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0561_),
    .Q_N(_3627_),
    .Q(rf_reg[609]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[60]_reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(rst_ni),
    .D(_0562_),
    .Q_N(_3626_),
    .Q(rf_reg[60]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[610]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0563_),
    .Q_N(_3625_),
    .Q(rf_reg[610]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[611]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0564_),
    .Q_N(_3624_),
    .Q(rf_reg[611]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[612]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0565_),
    .Q_N(_3623_),
    .Q(rf_reg[612]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[613]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0566_),
    .Q_N(_3622_),
    .Q(rf_reg[613]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[614]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0567_),
    .Q_N(_3621_),
    .Q(rf_reg[614]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[615]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0568_),
    .Q_N(_3620_),
    .Q(rf_reg[615]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[616]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0569_),
    .Q_N(_3619_),
    .Q(rf_reg[616]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[617]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0570_),
    .Q_N(_3618_),
    .Q(rf_reg[617]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[618]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0571_),
    .Q_N(_3617_),
    .Q(rf_reg[618]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[619]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0572_),
    .Q_N(_3616_),
    .Q(rf_reg[619]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[61]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0573_),
    .Q_N(_3615_),
    .Q(rf_reg[61]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[620]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0574_),
    .Q_N(_3614_),
    .Q(rf_reg[620]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[621]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0575_),
    .Q_N(_3613_),
    .Q(rf_reg[621]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[622]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0576_),
    .Q_N(_3612_),
    .Q(rf_reg[622]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[623]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0577_),
    .Q_N(_3611_),
    .Q(rf_reg[623]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[624]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0578_),
    .Q_N(_3610_),
    .Q(rf_reg[624]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[625]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0579_),
    .Q_N(_3609_),
    .Q(rf_reg[625]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[626]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0580_),
    .Q_N(_3608_),
    .Q(rf_reg[626]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[627]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0581_),
    .Q_N(_3607_),
    .Q(rf_reg[627]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[628]_reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(rst_ni),
    .D(_0582_),
    .Q_N(_3606_),
    .Q(rf_reg[628]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[629]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0583_),
    .Q_N(_3605_),
    .Q(rf_reg[629]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[62]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0584_),
    .Q_N(_3604_),
    .Q(rf_reg[62]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[630]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0585_),
    .Q_N(_3603_),
    .Q(rf_reg[630]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[631]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0586_),
    .Q_N(_3602_),
    .Q(rf_reg[631]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[632]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0587_),
    .Q_N(_3601_),
    .Q(rf_reg[632]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[633]_reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(rst_ni),
    .D(_0588_),
    .Q_N(_3600_),
    .Q(rf_reg[633]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[634]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0589_),
    .Q_N(_3599_),
    .Q(rf_reg[634]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[635]_reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(rst_ni),
    .D(_0590_),
    .Q_N(_3598_),
    .Q(rf_reg[635]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[636]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0591_),
    .Q_N(_3597_),
    .Q(rf_reg[636]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[637]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0592_),
    .Q_N(_3596_),
    .Q(rf_reg[637]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[638]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0593_),
    .Q_N(_3595_),
    .Q(rf_reg[638]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[639]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0594_),
    .Q_N(_3594_),
    .Q(rf_reg[639]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[63]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0595_),
    .Q_N(_3593_),
    .Q(rf_reg[63]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[640]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0596_),
    .Q_N(_3592_),
    .Q(rf_reg[640]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[641]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0597_),
    .Q_N(_3591_),
    .Q(rf_reg[641]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[642]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0598_),
    .Q_N(_3590_),
    .Q(rf_reg[642]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[643]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0599_),
    .Q_N(_3589_),
    .Q(rf_reg[643]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[644]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0600_),
    .Q_N(_3588_),
    .Q(rf_reg[644]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[645]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0601_),
    .Q_N(_3587_),
    .Q(rf_reg[645]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[646]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0602_),
    .Q_N(_3586_),
    .Q(rf_reg[646]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[647]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0603_),
    .Q_N(_3585_),
    .Q(rf_reg[647]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[648]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0604_),
    .Q_N(_3584_),
    .Q(rf_reg[648]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[649]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0605_),
    .Q_N(_3583_),
    .Q(rf_reg[649]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[64]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0606_),
    .Q_N(_3582_),
    .Q(rf_reg[64]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[650]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0607_),
    .Q_N(_3581_),
    .Q(rf_reg[650]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[651]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0608_),
    .Q_N(_3580_),
    .Q(rf_reg[651]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[652]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0609_),
    .Q_N(_3579_),
    .Q(rf_reg[652]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[653]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0610_),
    .Q_N(_3578_),
    .Q(rf_reg[653]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[654]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0611_),
    .Q_N(_3577_),
    .Q(rf_reg[654]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[655]_reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(rst_ni),
    .D(_0612_),
    .Q_N(_3576_),
    .Q(rf_reg[655]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[656]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0613_),
    .Q_N(_3575_),
    .Q(rf_reg[656]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[657]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0614_),
    .Q_N(_3574_),
    .Q(rf_reg[657]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[658]_reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(rst_ni),
    .D(_0615_),
    .Q_N(_3573_),
    .Q(rf_reg[658]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[659]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0616_),
    .Q_N(_3572_),
    .Q(rf_reg[659]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[65]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0617_),
    .Q_N(_3571_),
    .Q(rf_reg[65]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[660]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0618_),
    .Q_N(_3570_),
    .Q(rf_reg[660]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[661]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0619_),
    .Q_N(_3569_),
    .Q(rf_reg[661]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[662]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0620_),
    .Q_N(_3568_),
    .Q(rf_reg[662]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[663]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0621_),
    .Q_N(_3567_),
    .Q(rf_reg[663]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[664]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0622_),
    .Q_N(_3566_),
    .Q(rf_reg[664]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[665]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0623_),
    .Q_N(_3565_),
    .Q(rf_reg[665]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[666]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(_0624_),
    .Q_N(_3564_),
    .Q(rf_reg[666]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[667]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0625_),
    .Q_N(_3563_),
    .Q(rf_reg[667]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[668]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0626_),
    .Q_N(_3562_),
    .Q(rf_reg[668]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[669]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0627_),
    .Q_N(_3561_),
    .Q(rf_reg[669]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[66]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0628_),
    .Q_N(_3560_),
    .Q(rf_reg[66]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[670]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0629_),
    .Q_N(_3559_),
    .Q(rf_reg[670]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[671]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0630_),
    .Q_N(_3558_),
    .Q(rf_reg[671]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[672]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0631_),
    .Q_N(_3557_),
    .Q(rf_reg[672]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[673]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0632_),
    .Q_N(_3556_),
    .Q(rf_reg[673]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[674]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0633_),
    .Q_N(_3555_),
    .Q(rf_reg[674]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[675]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0634_),
    .Q_N(_3554_),
    .Q(rf_reg[675]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[676]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0635_),
    .Q_N(_3553_),
    .Q(rf_reg[676]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[677]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0636_),
    .Q_N(_3552_),
    .Q(rf_reg[677]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[678]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0637_),
    .Q_N(_3551_),
    .Q(rf_reg[678]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[679]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0638_),
    .Q_N(_3550_),
    .Q(rf_reg[679]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[67]_reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(rst_ni),
    .D(_0639_),
    .Q_N(_3549_),
    .Q(rf_reg[67]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[680]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0640_),
    .Q_N(_3548_),
    .Q(rf_reg[680]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[681]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0641_),
    .Q_N(_3547_),
    .Q(rf_reg[681]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[682]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0642_),
    .Q_N(_3546_),
    .Q(rf_reg[682]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[683]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0643_),
    .Q_N(_3545_),
    .Q(rf_reg[683]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[684]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0644_),
    .Q_N(_3544_),
    .Q(rf_reg[684]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[685]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0645_),
    .Q_N(_3543_),
    .Q(rf_reg[685]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[686]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0646_),
    .Q_N(_3542_),
    .Q(rf_reg[686]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[687]_reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(rst_ni),
    .D(_0647_),
    .Q_N(_3541_),
    .Q(rf_reg[687]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[688]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0648_),
    .Q_N(_3540_),
    .Q(rf_reg[688]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[689]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0649_),
    .Q_N(_3539_),
    .Q(rf_reg[689]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[68]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0650_),
    .Q_N(_3538_),
    .Q(rf_reg[68]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[690]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0651_),
    .Q_N(_3537_),
    .Q(rf_reg[690]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[691]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0652_),
    .Q_N(_3536_),
    .Q(rf_reg[691]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[692]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0653_),
    .Q_N(_3535_),
    .Q(rf_reg[692]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[693]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0654_),
    .Q_N(_3534_),
    .Q(rf_reg[693]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[694]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0655_),
    .Q_N(_3533_),
    .Q(rf_reg[694]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[695]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0656_),
    .Q_N(_3532_),
    .Q(rf_reg[695]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[696]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0657_),
    .Q_N(_3531_),
    .Q(rf_reg[696]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[697]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0658_),
    .Q_N(_3530_),
    .Q(rf_reg[697]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[698]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0659_),
    .Q_N(_3529_),
    .Q(rf_reg[698]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[699]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0660_),
    .Q_N(_3528_),
    .Q(rf_reg[699]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[69]_reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(rst_ni),
    .D(_0661_),
    .Q_N(_3527_),
    .Q(rf_reg[69]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[700]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0662_),
    .Q_N(_3526_),
    .Q(rf_reg[700]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[701]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0663_),
    .Q_N(_3525_),
    .Q(rf_reg[701]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[702]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0664_),
    .Q_N(_3524_),
    .Q(rf_reg[702]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[703]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0665_),
    .Q_N(_3523_),
    .Q(rf_reg[703]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[704]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0666_),
    .Q_N(_3522_),
    .Q(rf_reg[704]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[705]_reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(rst_ni),
    .D(_0667_),
    .Q_N(_3521_),
    .Q(rf_reg[705]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[706]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0668_),
    .Q_N(_3520_),
    .Q(rf_reg[706]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[707]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0669_),
    .Q_N(_3519_),
    .Q(rf_reg[707]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[708]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0670_),
    .Q_N(_3518_),
    .Q(rf_reg[708]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[709]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0671_),
    .Q_N(_3517_),
    .Q(rf_reg[709]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[70]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0672_),
    .Q_N(_3516_),
    .Q(rf_reg[70]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[710]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0673_),
    .Q_N(_3515_),
    .Q(rf_reg[710]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[711]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0674_),
    .Q_N(_3514_),
    .Q(rf_reg[711]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[712]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0675_),
    .Q_N(_3513_),
    .Q(rf_reg[712]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[713]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0676_),
    .Q_N(_3512_),
    .Q(rf_reg[713]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[714]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0677_),
    .Q_N(_3511_),
    .Q(rf_reg[714]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[715]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0678_),
    .Q_N(_3510_),
    .Q(rf_reg[715]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[716]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0679_),
    .Q_N(_3509_),
    .Q(rf_reg[716]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[717]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0680_),
    .Q_N(_3508_),
    .Q(rf_reg[717]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[718]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0681_),
    .Q_N(_3507_),
    .Q(rf_reg[718]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[719]_reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(rst_ni),
    .D(_0682_),
    .Q_N(_3506_),
    .Q(rf_reg[719]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[71]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0683_),
    .Q_N(_3505_),
    .Q(rf_reg[71]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[720]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0684_),
    .Q_N(_3504_),
    .Q(rf_reg[720]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[721]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0685_),
    .Q_N(_3503_),
    .Q(rf_reg[721]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[722]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0686_),
    .Q_N(_3502_),
    .Q(rf_reg[722]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[723]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0687_),
    .Q_N(_3501_),
    .Q(rf_reg[723]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[724]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0688_),
    .Q_N(_3500_),
    .Q(rf_reg[724]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[725]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0689_),
    .Q_N(_3499_),
    .Q(rf_reg[725]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[726]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0690_),
    .Q_N(_3498_),
    .Q(rf_reg[726]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[727]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0691_),
    .Q_N(_3497_),
    .Q(rf_reg[727]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[728]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0692_),
    .Q_N(_3496_),
    .Q(rf_reg[728]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[729]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0693_),
    .Q_N(_3495_),
    .Q(rf_reg[729]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[72]_reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(rst_ni),
    .D(_0694_),
    .Q_N(_3494_),
    .Q(rf_reg[72]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[730]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(_0695_),
    .Q_N(_3493_),
    .Q(rf_reg[730]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[731]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0696_),
    .Q_N(_3492_),
    .Q(rf_reg[731]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[732]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0697_),
    .Q_N(_3491_),
    .Q(rf_reg[732]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[733]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0698_),
    .Q_N(_3490_),
    .Q(rf_reg[733]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[734]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0699_),
    .Q_N(_3489_),
    .Q(rf_reg[734]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[735]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0700_),
    .Q_N(_3488_),
    .Q(rf_reg[735]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[736]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0701_),
    .Q_N(_3487_),
    .Q(rf_reg[736]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[737]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0702_),
    .Q_N(_3486_),
    .Q(rf_reg[737]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[738]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0703_),
    .Q_N(_3485_),
    .Q(rf_reg[738]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[739]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0704_),
    .Q_N(_3484_),
    .Q(rf_reg[739]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[73]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0705_),
    .Q_N(_3483_),
    .Q(rf_reg[73]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[740]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0706_),
    .Q_N(_3482_),
    .Q(rf_reg[740]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[741]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0707_),
    .Q_N(_3481_),
    .Q(rf_reg[741]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[742]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0708_),
    .Q_N(_3480_),
    .Q(rf_reg[742]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[743]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0709_),
    .Q_N(_3479_),
    .Q(rf_reg[743]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[744]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0710_),
    .Q_N(_3478_),
    .Q(rf_reg[744]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[745]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0711_),
    .Q_N(_3477_),
    .Q(rf_reg[745]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[746]_reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(rst_ni),
    .D(_0712_),
    .Q_N(_3476_),
    .Q(rf_reg[746]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[747]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0713_),
    .Q_N(_3475_),
    .Q(rf_reg[747]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[748]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0714_),
    .Q_N(_3474_),
    .Q(rf_reg[748]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[749]_reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(rst_ni),
    .D(_0715_),
    .Q_N(_3473_),
    .Q(rf_reg[749]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[74]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0716_),
    .Q_N(_3472_),
    .Q(rf_reg[74]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[750]_reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(rst_ni),
    .D(_0717_),
    .Q_N(_3471_),
    .Q(rf_reg[750]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[751]_reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(rst_ni),
    .D(_0718_),
    .Q_N(_3470_),
    .Q(rf_reg[751]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[752]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0719_),
    .Q_N(_3469_),
    .Q(rf_reg[752]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[753]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0720_),
    .Q_N(_3468_),
    .Q(rf_reg[753]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[754]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0721_),
    .Q_N(_3467_),
    .Q(rf_reg[754]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[755]_reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(rst_ni),
    .D(_0722_),
    .Q_N(_3466_),
    .Q(rf_reg[755]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[756]_reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(rst_ni),
    .D(_0723_),
    .Q_N(_3465_),
    .Q(rf_reg[756]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[757]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(_0724_),
    .Q_N(_3464_),
    .Q(rf_reg[757]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[758]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0725_),
    .Q_N(_3463_),
    .Q(rf_reg[758]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[759]_reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(rst_ni),
    .D(_0726_),
    .Q_N(_3462_),
    .Q(rf_reg[759]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[75]_reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(rst_ni),
    .D(_0727_),
    .Q_N(_3461_),
    .Q(rf_reg[75]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[760]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0728_),
    .Q_N(_3460_),
    .Q(rf_reg[760]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[761]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0729_),
    .Q_N(_3459_),
    .Q(rf_reg[761]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[762]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(_0730_),
    .Q_N(_3458_),
    .Q(rf_reg[762]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[763]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0731_),
    .Q_N(_3457_),
    .Q(rf_reg[763]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[764]_reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(rst_ni),
    .D(_0732_),
    .Q_N(_3456_),
    .Q(rf_reg[764]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[765]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0733_),
    .Q_N(_3455_),
    .Q(rf_reg[765]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[766]_reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(rst_ni),
    .D(_0734_),
    .Q_N(_3454_),
    .Q(rf_reg[766]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[767]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0735_),
    .Q_N(_3453_),
    .Q(rf_reg[767]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[768]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0736_),
    .Q_N(_3452_),
    .Q(rf_reg[768]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[769]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0737_),
    .Q_N(_3451_),
    .Q(rf_reg[769]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[76]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0738_),
    .Q_N(_3450_),
    .Q(rf_reg[76]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[770]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0739_),
    .Q_N(_3449_),
    .Q(rf_reg[770]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[771]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0740_),
    .Q_N(_3448_),
    .Q(rf_reg[771]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[772]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0741_),
    .Q_N(_3447_),
    .Q(rf_reg[772]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[773]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0742_),
    .Q_N(_3446_),
    .Q(rf_reg[773]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[774]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0743_),
    .Q_N(_3445_),
    .Q(rf_reg[774]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[775]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0744_),
    .Q_N(_3444_),
    .Q(rf_reg[775]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[776]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0745_),
    .Q_N(_3443_),
    .Q(rf_reg[776]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[777]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0746_),
    .Q_N(_3442_),
    .Q(rf_reg[777]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[778]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0747_),
    .Q_N(_3441_),
    .Q(rf_reg[778]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[779]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0748_),
    .Q_N(_3440_),
    .Q(rf_reg[779]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[77]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0749_),
    .Q_N(_3439_),
    .Q(rf_reg[77]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[780]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0750_),
    .Q_N(_3438_),
    .Q(rf_reg[780]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[781]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0751_),
    .Q_N(_3437_),
    .Q(rf_reg[781]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[782]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0752_),
    .Q_N(_3436_),
    .Q(rf_reg[782]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[783]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0753_),
    .Q_N(_3435_),
    .Q(rf_reg[783]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[784]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0754_),
    .Q_N(_3434_),
    .Q(rf_reg[784]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[785]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0755_),
    .Q_N(_3433_),
    .Q(rf_reg[785]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[786]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0756_),
    .Q_N(_3432_),
    .Q(rf_reg[786]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[787]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0757_),
    .Q_N(_3431_),
    .Q(rf_reg[787]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[788]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0758_),
    .Q_N(_3430_),
    .Q(rf_reg[788]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[789]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0759_),
    .Q_N(_3429_),
    .Q(rf_reg[789]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[78]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0760_),
    .Q_N(_3428_),
    .Q(rf_reg[78]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[790]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0761_),
    .Q_N(_3427_),
    .Q(rf_reg[790]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[791]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0762_),
    .Q_N(_3426_),
    .Q(rf_reg[791]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[792]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0763_),
    .Q_N(_3425_),
    .Q(rf_reg[792]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[793]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0764_),
    .Q_N(_3424_),
    .Q(rf_reg[793]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[794]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0765_),
    .Q_N(_3423_),
    .Q(rf_reg[794]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[795]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0766_),
    .Q_N(_3422_),
    .Q(rf_reg[795]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[796]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0767_),
    .Q_N(_3421_),
    .Q(rf_reg[796]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[797]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0768_),
    .Q_N(_3420_),
    .Q(rf_reg[797]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[798]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0769_),
    .Q_N(_3419_),
    .Q(rf_reg[798]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[799]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0770_),
    .Q_N(_3418_),
    .Q(rf_reg[799]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[79]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0771_),
    .Q_N(_3417_),
    .Q(rf_reg[79]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[800]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0772_),
    .Q_N(_3416_),
    .Q(rf_reg[800]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[801]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0773_),
    .Q_N(_3415_),
    .Q(rf_reg[801]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[802]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0774_),
    .Q_N(_3414_),
    .Q(rf_reg[802]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[803]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0775_),
    .Q_N(_3413_),
    .Q(rf_reg[803]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[804]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0776_),
    .Q_N(_3412_),
    .Q(rf_reg[804]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[805]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0777_),
    .Q_N(_3411_),
    .Q(rf_reg[805]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[806]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0778_),
    .Q_N(_3410_),
    .Q(rf_reg[806]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[807]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0779_),
    .Q_N(_3409_),
    .Q(rf_reg[807]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[808]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0780_),
    .Q_N(_3408_),
    .Q(rf_reg[808]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[809]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0781_),
    .Q_N(_3407_),
    .Q(rf_reg[809]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[80]_reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(rst_ni),
    .D(_0782_),
    .Q_N(_3406_),
    .Q(rf_reg[80]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[810]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0783_),
    .Q_N(_3405_),
    .Q(rf_reg[810]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[811]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0784_),
    .Q_N(_3404_),
    .Q(rf_reg[811]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[812]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0785_),
    .Q_N(_3403_),
    .Q(rf_reg[812]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[813]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0786_),
    .Q_N(_3402_),
    .Q(rf_reg[813]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[814]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0787_),
    .Q_N(_3401_),
    .Q(rf_reg[814]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[815]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0788_),
    .Q_N(_3400_),
    .Q(rf_reg[815]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[816]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0789_),
    .Q_N(_3399_),
    .Q(rf_reg[816]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[817]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0790_),
    .Q_N(_3398_),
    .Q(rf_reg[817]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[818]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0791_),
    .Q_N(_3397_),
    .Q(rf_reg[818]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[819]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0792_),
    .Q_N(_3396_),
    .Q(rf_reg[819]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[81]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0793_),
    .Q_N(_3395_),
    .Q(rf_reg[81]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[820]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0794_),
    .Q_N(_3394_),
    .Q(rf_reg[820]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[821]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0795_),
    .Q_N(_3393_),
    .Q(rf_reg[821]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[822]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(_0796_),
    .Q_N(_3392_),
    .Q(rf_reg[822]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[823]_reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(rst_ni),
    .D(_0797_),
    .Q_N(_3391_),
    .Q(rf_reg[823]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[824]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0798_),
    .Q_N(_3390_),
    .Q(rf_reg[824]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[825]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0799_),
    .Q_N(_3389_),
    .Q(rf_reg[825]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[826]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0800_),
    .Q_N(_3388_),
    .Q(rf_reg[826]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[827]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0801_),
    .Q_N(_3387_),
    .Q(rf_reg[827]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[828]_reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(rst_ni),
    .D(_0802_),
    .Q_N(_3386_),
    .Q(rf_reg[828]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[829]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0803_),
    .Q_N(_3385_),
    .Q(rf_reg[829]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[82]_reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(rst_ni),
    .D(_0804_),
    .Q_N(_3384_),
    .Q(rf_reg[82]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[830]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0805_),
    .Q_N(_3383_),
    .Q(rf_reg[830]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[831]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0806_),
    .Q_N(_3382_),
    .Q(rf_reg[831]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[832]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0807_),
    .Q_N(_3381_),
    .Q(rf_reg[832]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[833]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0808_),
    .Q_N(_3380_),
    .Q(rf_reg[833]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[834]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0809_),
    .Q_N(_3379_),
    .Q(rf_reg[834]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[835]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0810_),
    .Q_N(_3378_),
    .Q(rf_reg[835]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[836]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0811_),
    .Q_N(_3377_),
    .Q(rf_reg[836]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[837]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0812_),
    .Q_N(_3376_),
    .Q(rf_reg[837]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[838]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0813_),
    .Q_N(_3375_),
    .Q(rf_reg[838]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[839]_reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(rst_ni),
    .D(_0814_),
    .Q_N(_3374_),
    .Q(rf_reg[839]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[83]_reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(rst_ni),
    .D(_0815_),
    .Q_N(_3373_),
    .Q(rf_reg[83]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[840]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0816_),
    .Q_N(_3372_),
    .Q(rf_reg[840]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[841]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(_0817_),
    .Q_N(_3371_),
    .Q(rf_reg[841]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[842]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0818_),
    .Q_N(_3370_),
    .Q(rf_reg[842]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[843]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0819_),
    .Q_N(_3369_),
    .Q(rf_reg[843]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[844]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0820_),
    .Q_N(_3368_),
    .Q(rf_reg[844]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[845]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0821_),
    .Q_N(_3367_),
    .Q(rf_reg[845]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[846]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0822_),
    .Q_N(_3366_),
    .Q(rf_reg[846]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[847]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0823_),
    .Q_N(_3365_),
    .Q(rf_reg[847]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[848]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0824_),
    .Q_N(_3364_),
    .Q(rf_reg[848]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[849]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0825_),
    .Q_N(_3363_),
    .Q(rf_reg[849]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[84]_reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(rst_ni),
    .D(_0826_),
    .Q_N(_3362_),
    .Q(rf_reg[84]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[850]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0827_),
    .Q_N(_3361_),
    .Q(rf_reg[850]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[851]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0828_),
    .Q_N(_3360_),
    .Q(rf_reg[851]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[852]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0829_),
    .Q_N(_3359_),
    .Q(rf_reg[852]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[853]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0830_),
    .Q_N(_3358_),
    .Q(rf_reg[853]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[854]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0831_),
    .Q_N(_3357_),
    .Q(rf_reg[854]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[855]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0832_),
    .Q_N(_3356_),
    .Q(rf_reg[855]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[856]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0833_),
    .Q_N(_3355_),
    .Q(rf_reg[856]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[857]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0834_),
    .Q_N(_3354_),
    .Q(rf_reg[857]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[858]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0835_),
    .Q_N(_3353_),
    .Q(rf_reg[858]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[859]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0836_),
    .Q_N(_3352_),
    .Q(rf_reg[859]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[85]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0837_),
    .Q_N(_3351_),
    .Q(rf_reg[85]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[860]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0838_),
    .Q_N(_3350_),
    .Q(rf_reg[860]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[861]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0839_),
    .Q_N(_3349_),
    .Q(rf_reg[861]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[862]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0840_),
    .Q_N(_3348_),
    .Q(rf_reg[862]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[863]_reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(rst_ni),
    .D(_0841_),
    .Q_N(_3347_),
    .Q(rf_reg[863]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[864]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0842_),
    .Q_N(_3346_),
    .Q(rf_reg[864]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[865]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0843_),
    .Q_N(_3345_),
    .Q(rf_reg[865]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[866]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0844_),
    .Q_N(_3344_),
    .Q(rf_reg[866]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[867]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0845_),
    .Q_N(_3343_),
    .Q(rf_reg[867]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[868]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0846_),
    .Q_N(_3342_),
    .Q(rf_reg[868]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[869]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0847_),
    .Q_N(_3341_),
    .Q(rf_reg[869]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[86]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0848_),
    .Q_N(_3340_),
    .Q(rf_reg[86]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[870]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0849_),
    .Q_N(_3339_),
    .Q(rf_reg[870]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[871]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0850_),
    .Q_N(_3338_),
    .Q(rf_reg[871]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[872]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0851_),
    .Q_N(_3337_),
    .Q(rf_reg[872]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[873]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0852_),
    .Q_N(_3336_),
    .Q(rf_reg[873]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[874]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(_0853_),
    .Q_N(_3335_),
    .Q(rf_reg[874]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[875]_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(rst_ni),
    .D(_0854_),
    .Q_N(_3334_),
    .Q(rf_reg[875]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[876]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0855_),
    .Q_N(_3333_),
    .Q(rf_reg[876]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[877]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0856_),
    .Q_N(_3332_),
    .Q(rf_reg[877]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[878]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0857_),
    .Q_N(_3331_),
    .Q(rf_reg[878]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[879]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0858_),
    .Q_N(_3330_),
    .Q(rf_reg[879]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[87]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0859_),
    .Q_N(_3329_),
    .Q(rf_reg[87]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[880]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0860_),
    .Q_N(_3328_),
    .Q(rf_reg[880]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[881]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0861_),
    .Q_N(_3327_),
    .Q(rf_reg[881]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[882]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0862_),
    .Q_N(_3326_),
    .Q(rf_reg[882]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[883]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0863_),
    .Q_N(_3325_),
    .Q(rf_reg[883]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[884]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0864_),
    .Q_N(_3324_),
    .Q(rf_reg[884]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[885]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0865_),
    .Q_N(_3323_),
    .Q(rf_reg[885]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[886]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0866_),
    .Q_N(_3322_),
    .Q(rf_reg[886]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[887]_reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(rst_ni),
    .D(_0867_),
    .Q_N(_3321_),
    .Q(rf_reg[887]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[888]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0868_),
    .Q_N(_3320_),
    .Q(rf_reg[888]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[889]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0869_),
    .Q_N(_3319_),
    .Q(rf_reg[889]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[88]_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(rst_ni),
    .D(_0870_),
    .Q_N(_3318_),
    .Q(rf_reg[88]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[890]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0871_),
    .Q_N(_3317_),
    .Q(rf_reg[890]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[891]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0872_),
    .Q_N(_3316_),
    .Q(rf_reg[891]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[892]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0873_),
    .Q_N(_3315_),
    .Q(rf_reg[892]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[893]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0874_),
    .Q_N(_3314_),
    .Q(rf_reg[893]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[894]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0875_),
    .Q_N(_3313_),
    .Q(rf_reg[894]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[895]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(_0876_),
    .Q_N(_3312_),
    .Q(rf_reg[895]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[896]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0877_),
    .Q_N(_3311_),
    .Q(rf_reg[896]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[897]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0878_),
    .Q_N(_3310_),
    .Q(rf_reg[897]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[898]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0879_),
    .Q_N(_3309_),
    .Q(rf_reg[898]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[899]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0880_),
    .Q_N(_3308_),
    .Q(rf_reg[899]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[89]_reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(rst_ni),
    .D(_0881_),
    .Q_N(_3307_),
    .Q(rf_reg[89]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[900]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0882_),
    .Q_N(_3306_),
    .Q(rf_reg[900]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[901]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0883_),
    .Q_N(_3305_),
    .Q(rf_reg[901]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[902]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0884_),
    .Q_N(_3304_),
    .Q(rf_reg[902]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[903]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0885_),
    .Q_N(_3303_),
    .Q(rf_reg[903]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[904]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0886_),
    .Q_N(_3302_),
    .Q(rf_reg[904]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[905]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(_0887_),
    .Q_N(_3301_),
    .Q(rf_reg[905]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[906]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0888_),
    .Q_N(_3300_),
    .Q(rf_reg[906]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[907]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0889_),
    .Q_N(_3299_),
    .Q(rf_reg[907]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[908]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0890_),
    .Q_N(_3298_),
    .Q(rf_reg[908]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[909]_reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(rst_ni),
    .D(_0891_),
    .Q_N(_3297_),
    .Q(rf_reg[909]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[90]_reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(rst_ni),
    .D(_0892_),
    .Q_N(_3296_),
    .Q(rf_reg[90]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[910]_reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(rst_ni),
    .D(_0893_),
    .Q_N(_3295_),
    .Q(rf_reg[910]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[911]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0894_),
    .Q_N(_3294_),
    .Q(rf_reg[911]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[912]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0895_),
    .Q_N(_3293_),
    .Q(rf_reg[912]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[913]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0896_),
    .Q_N(_3292_),
    .Q(rf_reg[913]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[914]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0897_),
    .Q_N(_3291_),
    .Q(rf_reg[914]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[915]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0898_),
    .Q_N(_3290_),
    .Q(rf_reg[915]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[916]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0899_),
    .Q_N(_3289_),
    .Q(rf_reg[916]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[917]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0900_),
    .Q_N(_3288_),
    .Q(rf_reg[917]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[918]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0901_),
    .Q_N(_3287_),
    .Q(rf_reg[918]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[919]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0902_),
    .Q_N(_3286_),
    .Q(rf_reg[919]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[91]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0903_),
    .Q_N(_3285_),
    .Q(rf_reg[91]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[920]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0904_),
    .Q_N(_3284_),
    .Q(rf_reg[920]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[921]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0905_),
    .Q_N(_3283_),
    .Q(rf_reg[921]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[922]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0906_),
    .Q_N(_3282_),
    .Q(rf_reg[922]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[923]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0907_),
    .Q_N(_3281_),
    .Q(rf_reg[923]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[924]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0908_),
    .Q_N(_3280_),
    .Q(rf_reg[924]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[925]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0909_),
    .Q_N(_3279_),
    .Q(rf_reg[925]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[926]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0910_),
    .Q_N(_3278_),
    .Q(rf_reg[926]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[927]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0911_),
    .Q_N(_3277_),
    .Q(rf_reg[927]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[928]_reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(rst_ni),
    .D(_0912_),
    .Q_N(_3276_),
    .Q(rf_reg[928]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[929]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0913_),
    .Q_N(_3275_),
    .Q(rf_reg[929]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[92]_reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(rst_ni),
    .D(_0914_),
    .Q_N(_3274_),
    .Q(rf_reg[92]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[930]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0915_),
    .Q_N(_3273_),
    .Q(rf_reg[930]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[931]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0916_),
    .Q_N(_3272_),
    .Q(rf_reg[931]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[932]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0917_),
    .Q_N(_3271_),
    .Q(rf_reg[932]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[933]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0918_),
    .Q_N(_3270_),
    .Q(rf_reg[933]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[934]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0919_),
    .Q_N(_3269_),
    .Q(rf_reg[934]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[935]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0920_),
    .Q_N(_3268_),
    .Q(rf_reg[935]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[936]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0921_),
    .Q_N(_3267_),
    .Q(rf_reg[936]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[937]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(_0922_),
    .Q_N(_3266_),
    .Q(rf_reg[937]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[938]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0923_),
    .Q_N(_3265_),
    .Q(rf_reg[938]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[939]_reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(rst_ni),
    .D(_0924_),
    .Q_N(_3264_),
    .Q(rf_reg[939]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[93]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0925_),
    .Q_N(_3263_),
    .Q(rf_reg[93]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[940]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0926_),
    .Q_N(_3262_),
    .Q(rf_reg[940]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[941]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0927_),
    .Q_N(_3261_),
    .Q(rf_reg[941]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[942]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0928_),
    .Q_N(_3260_),
    .Q(rf_reg[942]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[943]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0929_),
    .Q_N(_3259_),
    .Q(rf_reg[943]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[944]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0930_),
    .Q_N(_3258_),
    .Q(rf_reg[944]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[945]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(_0931_),
    .Q_N(_3257_),
    .Q(rf_reg[945]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[946]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0932_),
    .Q_N(_3256_),
    .Q(rf_reg[946]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[947]_reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(rst_ni),
    .D(_0933_),
    .Q_N(_3255_),
    .Q(rf_reg[947]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[948]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0934_),
    .Q_N(_3254_),
    .Q(rf_reg[948]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[949]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(_0935_),
    .Q_N(_3253_),
    .Q(rf_reg[949]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[94]_reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(rst_ni),
    .D(_0936_),
    .Q_N(_3252_),
    .Q(rf_reg[94]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[950]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0937_),
    .Q_N(_3251_),
    .Q(rf_reg[950]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[951]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0938_),
    .Q_N(_3250_),
    .Q(rf_reg[951]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[952]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0939_),
    .Q_N(_3249_),
    .Q(rf_reg[952]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[953]_reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(rst_ni),
    .D(_0940_),
    .Q_N(_3248_),
    .Q(rf_reg[953]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[954]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0941_),
    .Q_N(_3247_),
    .Q(rf_reg[954]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[955]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0942_),
    .Q_N(_3246_),
    .Q(rf_reg[955]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[956]_reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(rst_ni),
    .D(_0943_),
    .Q_N(_3245_),
    .Q(rf_reg[956]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[957]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0944_),
    .Q_N(_3244_),
    .Q(rf_reg[957]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[958]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0945_),
    .Q_N(_3243_),
    .Q(rf_reg[958]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[959]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0946_),
    .Q_N(_3242_),
    .Q(rf_reg[959]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[95]_reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(rst_ni),
    .D(_0947_),
    .Q_N(_3241_),
    .Q(rf_reg[95]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[960]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0948_),
    .Q_N(_3240_),
    .Q(rf_reg[960]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[961]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0949_),
    .Q_N(_3239_),
    .Q(rf_reg[961]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[962]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0950_),
    .Q_N(_3238_),
    .Q(rf_reg[962]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[963]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0951_),
    .Q_N(_3237_),
    .Q(rf_reg[963]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[964]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0952_),
    .Q_N(_3236_),
    .Q(rf_reg[964]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[965]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0953_),
    .Q_N(_3235_),
    .Q(rf_reg[965]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[966]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0954_),
    .Q_N(_3234_),
    .Q(rf_reg[966]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[967]_reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(rst_ni),
    .D(_0955_),
    .Q_N(_3233_),
    .Q(rf_reg[967]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[968]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0956_),
    .Q_N(_3232_),
    .Q(rf_reg[968]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[969]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(_0957_),
    .Q_N(_3231_),
    .Q(rf_reg[969]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[96]_reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(rst_ni),
    .D(_0958_),
    .Q_N(_3230_),
    .Q(rf_reg[96]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[970]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0959_),
    .Q_N(_3229_),
    .Q(rf_reg[970]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[971]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0960_),
    .Q_N(_3228_),
    .Q(rf_reg[971]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[972]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0961_),
    .Q_N(_3227_),
    .Q(rf_reg[972]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[973]_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(rst_ni),
    .D(_0962_),
    .Q_N(_3226_),
    .Q(rf_reg[973]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[974]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0963_),
    .Q_N(_3225_),
    .Q(rf_reg[974]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[975]_reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(rst_ni),
    .D(_0964_),
    .Q_N(_3224_),
    .Q(rf_reg[975]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[976]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0965_),
    .Q_N(_3223_),
    .Q(rf_reg[976]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[977]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0966_),
    .Q_N(_3222_),
    .Q(rf_reg[977]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[978]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0967_),
    .Q_N(_3221_),
    .Q(rf_reg[978]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[979]_reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(rst_ni),
    .D(_0968_),
    .Q_N(_3220_),
    .Q(rf_reg[979]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[97]_reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(rst_ni),
    .D(_0969_),
    .Q_N(_3219_),
    .Q(rf_reg[97]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[980]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0970_),
    .Q_N(_3218_),
    .Q(rf_reg[980]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[981]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0971_),
    .Q_N(_3217_),
    .Q(rf_reg[981]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[982]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0972_),
    .Q_N(_3216_),
    .Q(rf_reg[982]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[983]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0973_),
    .Q_N(_3215_),
    .Q(rf_reg[983]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[984]_reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(rst_ni),
    .D(_0974_),
    .Q_N(_3214_),
    .Q(rf_reg[984]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[985]_reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(rst_ni),
    .D(_0975_),
    .Q_N(_3213_),
    .Q(rf_reg[985]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[986]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0976_),
    .Q_N(_3212_),
    .Q(rf_reg[986]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[987]_reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(rst_ni),
    .D(_0977_),
    .Q_N(_3211_),
    .Q(rf_reg[987]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[988]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0978_),
    .Q_N(_3210_),
    .Q(rf_reg[988]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[989]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0979_),
    .Q_N(_3209_),
    .Q(rf_reg[989]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[98]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0980_),
    .Q_N(_3208_),
    .Q(rf_reg[98]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[990]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(_0981_),
    .Q_N(_3207_),
    .Q(rf_reg[990]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[991]_reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(rst_ni),
    .D(_0982_),
    .Q_N(_3206_),
    .Q(rf_reg[991]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[992]_reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(rst_ni),
    .D(_0983_),
    .Q_N(_3205_),
    .Q(rf_reg[992]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[993]_reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(rst_ni),
    .D(_0984_),
    .Q_N(_3204_),
    .Q(rf_reg[993]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[994]_reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(rst_ni),
    .D(_0985_),
    .Q_N(_3203_),
    .Q(rf_reg[994]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[995]_reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(rst_ni),
    .D(_0986_),
    .Q_N(_3202_),
    .Q(rf_reg[995]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[996]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0987_),
    .Q_N(_3201_),
    .Q(rf_reg[996]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[997]_reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(rst_ni),
    .D(_0988_),
    .Q_N(_3200_),
    .Q(rf_reg[997]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[998]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(_0989_),
    .Q_N(_3199_),
    .Q(rf_reg[998]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[999]_reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(rst_ni),
    .D(_0990_),
    .Q_N(_3198_),
    .Q(rf_reg[999]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \rf_reg[99]_reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(rst_ni),
    .D(_0991_),
    .Q_N(_3197_),
    .Q(rf_reg[99]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_124_clk_i (.X(clknet_leaf_124_clk_i),
    .A(clknet_5_4__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_125_clk_i (.X(clknet_leaf_125_clk_i),
    .A(clknet_5_4__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_126_clk_i (.X(clknet_leaf_126_clk_i),
    .A(clknet_5_4__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_127_clk_i (.X(clknet_leaf_127_clk_i),
    .A(clknet_5_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_128_clk_i (.X(clknet_leaf_128_clk_i),
    .A(clknet_5_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_129_clk_i (.X(clknet_leaf_129_clk_i),
    .A(clknet_5_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_leaf_130_clk_i (.X(clknet_leaf_130_clk_i),
    .A(clknet_5_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_0_0_clk_i (.X(clknet_4_0_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_1_0_clk_i (.X(clknet_4_1_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_2_0_clk_i (.X(clknet_4_2_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_3_0_clk_i (.X(clknet_4_3_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_4_0_clk_i (.X(clknet_4_4_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_5_0_clk_i (.X(clknet_4_5_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_6_0_clk_i (.X(clknet_4_6_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_7_0_clk_i (.X(clknet_4_7_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_8_0_clk_i (.X(clknet_4_8_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_9_0_clk_i (.X(clknet_4_9_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_10_0_clk_i (.X(clknet_4_10_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_11_0_clk_i (.X(clknet_4_11_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_12_0_clk_i (.X(clknet_4_12_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_13_0_clk_i (.X(clknet_4_13_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_14_0_clk_i (.X(clknet_4_14_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_4_15_0_clk_i (.X(clknet_4_15_0_clk_i),
    .A(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_0__f_clk_i (.A(clknet_4_0_0_clk_i),
    .X(clknet_5_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_1__f_clk_i (.A(clknet_4_0_0_clk_i),
    .X(clknet_5_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_2__f_clk_i (.A(clknet_4_1_0_clk_i),
    .X(clknet_5_2__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_3__f_clk_i (.A(clknet_4_1_0_clk_i),
    .X(clknet_5_3__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_4__f_clk_i (.A(clknet_4_2_0_clk_i),
    .X(clknet_5_4__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_5__f_clk_i (.A(clknet_4_2_0_clk_i),
    .X(clknet_5_5__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_6__f_clk_i (.A(clknet_4_3_0_clk_i),
    .X(clknet_5_6__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_7__f_clk_i (.A(clknet_4_3_0_clk_i),
    .X(clknet_5_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_8__f_clk_i (.A(clknet_4_4_0_clk_i),
    .X(clknet_5_8__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_9__f_clk_i (.A(clknet_4_4_0_clk_i),
    .X(clknet_5_9__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_10__f_clk_i (.A(clknet_4_5_0_clk_i),
    .X(clknet_5_10__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_11__f_clk_i (.A(clknet_4_5_0_clk_i),
    .X(clknet_5_11__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_12__f_clk_i (.A(clknet_4_6_0_clk_i),
    .X(clknet_5_12__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_13__f_clk_i (.A(clknet_4_6_0_clk_i),
    .X(clknet_5_13__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_14__f_clk_i (.A(clknet_4_7_0_clk_i),
    .X(clknet_5_14__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_15__f_clk_i (.A(clknet_4_7_0_clk_i),
    .X(clknet_5_15__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_16__f_clk_i (.A(clknet_4_8_0_clk_i),
    .X(clknet_5_16__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_17__f_clk_i (.A(clknet_4_8_0_clk_i),
    .X(clknet_5_17__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_18__f_clk_i (.A(clknet_4_9_0_clk_i),
    .X(clknet_5_18__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_19__f_clk_i (.A(clknet_4_9_0_clk_i),
    .X(clknet_5_19__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_20__f_clk_i (.A(clknet_4_10_0_clk_i),
    .X(clknet_5_20__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_21__f_clk_i (.A(clknet_4_10_0_clk_i),
    .X(clknet_5_21__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_22__f_clk_i (.A(clknet_4_11_0_clk_i),
    .X(clknet_5_22__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_23__f_clk_i (.A(clknet_4_11_0_clk_i),
    .X(clknet_5_23__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_24__f_clk_i (.A(clknet_4_12_0_clk_i),
    .X(clknet_5_24__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_25__f_clk_i (.A(clknet_4_12_0_clk_i),
    .X(clknet_5_25__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_26__f_clk_i (.A(clknet_4_13_0_clk_i),
    .X(clknet_5_26__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_27__f_clk_i (.A(clknet_4_13_0_clk_i),
    .X(clknet_5_27__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_28__f_clk_i (.A(clknet_4_14_0_clk_i),
    .X(clknet_5_28__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_29__f_clk_i (.A(clknet_4_14_0_clk_i),
    .X(clknet_5_29__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_30__f_clk_i (.A(clknet_4_15_0_clk_i),
    .X(clknet_5_30__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_5_31__f_clk_i (.A(clknet_4_15_0_clk_i),
    .X(clknet_5_31__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload0 (.A(clknet_5_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload1 (.A(clknet_5_9__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkload2 (.A(clknet_5_17__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_127_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload5 (.VDD(VDD),
    .A(clknet_leaf_8_clk_i),
    .VSS(VSS));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_11_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload7 (.VDD(VDD),
    .A(clknet_leaf_12_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload8 (.VDD(VDD),
    .A(clknet_leaf_125_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_126_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload10 (.VDD(VDD),
    .A(clknet_leaf_121_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload11 (.VDD(VDD),
    .A(clknet_leaf_123_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload12 (.VDD(VDD),
    .A(clknet_leaf_13_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload13 (.VDD(VDD),
    .A(clknet_leaf_118_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_115_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_26_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload16 (.VDD(VDD),
    .A(clknet_leaf_27_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload17 (.VDD(VDD),
    .A(clknet_leaf_31_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_33_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload19 (.VDD(VDD),
    .A(clknet_leaf_47_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload20 (.VDD(VDD),
    .A(clknet_leaf_46_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload21 (.VDD(VDD),
    .A(clknet_leaf_37_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload22 (.VDD(VDD),
    .A(clknet_leaf_39_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload23 (.VDD(VDD),
    .A(clknet_leaf_106_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_102_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_103_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload26 (.VDD(VDD),
    .A(clknet_leaf_113_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload27 (.VDD(VDD),
    .A(clknet_leaf_84_clk_i),
    .VSS(VSS));
 sg13g2_buf_8 clkload28 (.A(clknet_leaf_111_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload29 (.A(clknet_leaf_94_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload30 (.A(clknet_leaf_101_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload31 (.VDD(VDD),
    .A(clknet_leaf_96_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload32 (.VDD(VDD),
    .A(clknet_leaf_97_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload33 (.VDD(VDD),
    .A(clknet_leaf_90_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload34 (.VDD(VDD),
    .A(clknet_leaf_78_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload35 (.VDD(VDD),
    .A(clknet_leaf_79_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_63_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload37 (.A(clknet_leaf_65_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload38 (.VDD(VDD),
    .A(clknet_leaf_66_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_67_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd3_1 hold316 (.A(wdata_a_i[27]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold317 (.A(wdata_a_i[11]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold318 (.A(wdata_a_i[18]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold319 (.A(wdata_a_i[30]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold320 (.A(wdata_a_i[16]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold321 (.A(wdata_a_i[14]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold322 (.A(wdata_a_i[12]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold323 (.A(wdata_a_i[31]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold324 (.A(wdata_a_i[23]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold325 (.A(wdata_a_i[19]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold326 (.A(wdata_a_i[6]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold327 (.A(wdata_a_i[10]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold328 (.A(wdata_a_i[0]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold329 (.A(wdata_a_i[1]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold330 (.A(wdata_a_i[17]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold331 (.A(wdata_a_i[3]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold332 (.A(wdata_a_i[15]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold333 (.A(wdata_a_i[25]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold334 (.A(wdata_a_i[21]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold335 (.A(wdata_a_i[29]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold336 (.A(wdata_a_i[24]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold337 (.A(wdata_a_i[4]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold338 (.A(wdata_a_i[22]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold339 (.A(wdata_a_i[28]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold340 (.A(wdata_a_i[7]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold341 (.A(wdata_a_i[8]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold342 (.A(wdata_a_i[5]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold343 (.A(wdata_a_i[26]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold344 (.A(wdata_a_i[20]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold345 (.A(wdata_a_i[13]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold346 (.A(wdata_a_i[2]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold347 (.A(wdata_a_i[9]),
    .VDD(VDD),
    .VSS(VSS),
    .X(net347));
 sg13g2_antennanp ANTENNA_1 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[13]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[17]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[20]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[20]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[21]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[22]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[26]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[27]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[28]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[29]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[2]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[2]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[5]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[9]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[13]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[20]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[20]));
 sg13g2_antennanp ANTENNA_18 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[22]));
 sg13g2_antennanp ANTENNA_19 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[26]));
 sg13g2_antennanp ANTENNA_20 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[27]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[28]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[2]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[5]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[9]));
 sg13g2_antennanp ANTENNA_25 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[13]));
 sg13g2_antennanp ANTENNA_26 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[13]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[20]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[20]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[22]));
 sg13g2_antennanp ANTENNA_30 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[26]));
 sg13g2_antennanp ANTENNA_31 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[27]));
 sg13g2_antennanp ANTENNA_32 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[28]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[2]));
 sg13g2_antennanp ANTENNA_34 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[5]));
 sg13g2_antennanp ANTENNA_35 (.VDD(VDD),
    .VSS(VSS),
    .A(wdata_a_i[9]));
endmodule
