VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO cve2_register_file_ff
  FOREIGN cve2_register_file_ff 0 0 ;
  CLASS BLOCK ;
  SIZE 404.64 BY 410 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
  END VSS
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  286.94 409.28 287.14 410 ;
    END
  END clk_i
  PIN raddr_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  131.42 409.28 131.62 410 ;
    END
  END raddr_a_i[0]
  PIN raddr_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  141.5 409.28 141.7 410 ;
    END
  END raddr_a_i[1]
  PIN raddr_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  207.74 409.28 207.94 410 ;
    END
  END raddr_a_i[2]
  PIN raddr_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  127.1 409.28 127.3 410 ;
    END
  END raddr_a_i[3]
  PIN raddr_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  203.42 409.28 203.62 410 ;
    END
  END raddr_a_i[4]
  PIN raddr_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  210.62 409.28 210.82 410 ;
    END
  END raddr_b_i[0]
  PIN raddr_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  212.06 409.28 212.26 410 ;
    END
  END raddr_b_i[1]
  PIN raddr_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  213.5 409.28 213.7 410 ;
    END
  END raddr_b_i[2]
  PIN raddr_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  161.66 409.28 161.86 410 ;
    END
  END raddr_b_i[3]
  PIN raddr_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  214.94 409.28 215.14 410 ;
    END
  END raddr_b_i[4]
  PIN rdata_a_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  216.38 409.28 216.58 410 ;
    END
  END rdata_a_o[0]
  PIN rdata_a_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  217.82 409.28 218.02 410 ;
    END
  END rdata_a_o[10]
  PIN rdata_a_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  200.54 409.28 200.74 410 ;
    END
  END rdata_a_o[11]
  PIN rdata_a_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  160.22 409.28 160.42 410 ;
    END
  END rdata_a_o[12]
  PIN rdata_a_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  220.7 409.28 220.9 410 ;
    END
  END rdata_a_o[13]
  PIN rdata_a_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  140.06 409.28 140.26 410 ;
    END
  END rdata_a_o[14]
  PIN rdata_a_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  199.1 409.28 199.3 410 ;
    END
  END rdata_a_o[15]
  PIN rdata_a_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  181.82 409.28 182.02 410 ;
    END
  END rdata_a_o[16]
  PIN rdata_a_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  124.22 409.28 124.42 410 ;
    END
  END rdata_a_o[17]
  PIN rdata_a_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  226.46 409.28 226.66 410 ;
    END
  END rdata_a_o[18]
  PIN rdata_a_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  197.66 409.28 197.86 410 ;
    END
  END rdata_a_o[19]
  PIN rdata_a_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  227.9 409.28 228.1 410 ;
    END
  END rdata_a_o[1]
  PIN rdata_a_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  229.34 409.28 229.54 410 ;
    END
  END rdata_a_o[20]
  PIN rdata_a_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  157.34 409.28 157.54 410 ;
    END
  END rdata_a_o[21]
  PIN rdata_a_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  129.98 409.28 130.18 410 ;
    END
  END rdata_a_o[22]
  PIN rdata_a_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  232.22 409.28 232.42 410 ;
    END
  END rdata_a_o[23]
  PIN rdata_a_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  233.66 409.28 233.86 410 ;
    END
  END rdata_a_o[24]
  PIN rdata_a_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  138.62 409.28 138.82 410 ;
    END
  END rdata_a_o[25]
  PIN rdata_a_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  155.9 409.28 156.1 410 ;
    END
  END rdata_a_o[26]
  PIN rdata_a_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  236.54 409.28 236.74 410 ;
    END
  END rdata_a_o[27]
  PIN rdata_a_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  237.98 409.28 238.18 410 ;
    END
  END rdata_a_o[28]
  PIN rdata_a_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  154.46 409.28 154.66 410 ;
    END
  END rdata_a_o[29]
  PIN rdata_a_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  193.34 409.28 193.54 410 ;
    END
  END rdata_a_o[2]
  PIN rdata_a_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  151.58 409.28 151.78 410 ;
    END
  END rdata_a_o[30]
  PIN rdata_a_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  242.3 409.28 242.5 410 ;
    END
  END rdata_a_o[31]
  PIN rdata_a_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  243.74 409.28 243.94 410 ;
    END
  END rdata_a_o[3]
  PIN rdata_a_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  191.9 409.28 192.1 410 ;
    END
  END rdata_a_o[4]
  PIN rdata_a_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  245.18 409.28 245.38 410 ;
    END
  END rdata_a_o[5]
  PIN rdata_a_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  153.02 409.28 153.22 410 ;
    END
  END rdata_a_o[6]
  PIN rdata_a_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  248.06 409.28 248.26 410 ;
    END
  END rdata_a_o[7]
  PIN rdata_a_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  190.46 409.28 190.66 410 ;
    END
  END rdata_a_o[8]
  PIN rdata_a_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  187.58 409.28 187.78 410 ;
    END
  END rdata_a_o[9]
  PIN rdata_b_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  235.1 409.28 235.3 410 ;
    END
  END rdata_b_o[0]
  PIN rdata_b_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  137.18 409.28 137.38 410 ;
    END
  END rdata_b_o[10]
  PIN rdata_b_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  189.02 409.28 189.22 410 ;
    END
  END rdata_b_o[11]
  PIN rdata_b_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  204.86 409.28 205.06 410 ;
    END
  END rdata_b_o[12]
  PIN rdata_b_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  255.26 409.28 255.46 410 ;
    END
  END rdata_b_o[13]
  PIN rdata_b_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  256.7 409.28 256.9 410 ;
    END
  END rdata_b_o[14]
  PIN rdata_b_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  178.94 409.28 179.14 410 ;
    END
  END rdata_b_o[15]
  PIN rdata_b_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  222.14 409.28 222.34 410 ;
    END
  END rdata_b_o[16]
  PIN rdata_b_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  239.42 409.28 239.62 410 ;
    END
  END rdata_b_o[17]
  PIN rdata_b_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  150.14 409.28 150.34 410 ;
    END
  END rdata_b_o[18]
  PIN rdata_b_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  186.14 409.28 186.34 410 ;
    END
  END rdata_b_o[19]
  PIN rdata_b_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  183.26 409.28 183.46 410 ;
    END
  END rdata_b_o[1]
  PIN rdata_b_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  262.46 409.28 262.66 410 ;
    END
  END rdata_b_o[20]
  PIN rdata_b_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  135.74 409.28 135.94 410 ;
    END
  END rdata_b_o[21]
  PIN rdata_b_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  184.7 409.28 184.9 410 ;
    END
  END rdata_b_o[22]
  PIN rdata_b_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  206.3 409.28 206.5 410 ;
    END
  END rdata_b_o[23]
  PIN rdata_b_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  246.62 409.28 246.82 410 ;
    END
  END rdata_b_o[24]
  PIN rdata_b_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  265.34 409.28 265.54 410 ;
    END
  END rdata_b_o[25]
  PIN rdata_b_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  174.62 409.28 174.82 410 ;
    END
  END rdata_b_o[26]
  PIN rdata_b_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  148.7 409.28 148.9 410 ;
    END
  END rdata_b_o[27]
  PIN rdata_b_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  266.78 409.28 266.98 410 ;
    END
  END rdata_b_o[28]
  PIN rdata_b_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  171.74 409.28 171.94 410 ;
    END
  END rdata_b_o[29]
  PIN rdata_b_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  128.54 409.28 128.74 410 ;
    END
  END rdata_b_o[2]
  PIN rdata_b_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  230.78 409.28 230.98 410 ;
    END
  END rdata_b_o[30]
  PIN rdata_b_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  134.3 409.28 134.5 410 ;
    END
  END rdata_b_o[31]
  PIN rdata_b_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  225.02 409.28 225.22 410 ;
    END
  END rdata_b_o[3]
  PIN rdata_b_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  180.38 409.28 180.58 410 ;
    END
  END rdata_b_o[4]
  PIN rdata_b_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  269.66 409.28 269.86 410 ;
    END
  END rdata_b_o[5]
  PIN rdata_b_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  219.26 409.28 219.46 410 ;
    END
  END rdata_b_o[6]
  PIN rdata_b_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  253.82 409.28 254.02 410 ;
    END
  END rdata_b_o[7]
  PIN rdata_b_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  147.26 409.28 147.46 410 ;
    END
  END rdata_b_o[8]
  PIN rdata_b_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  125.66 409.28 125.86 410 ;
    END
  END rdata_b_o[9]
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  209.18 409.28 209.38 410 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1.82 0 2.02 0.72 ;
    END
  END test_en_i
  PIN waddr_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  263.9 409.28 264.1 410 ;
    END
  END waddr_a_i[0]
  PIN waddr_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  177.5 409.28 177.7 410 ;
    END
  END waddr_a_i[1]
  PIN waddr_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  196.22 409.28 196.42 410 ;
    END
  END waddr_a_i[2]
  PIN waddr_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  273.98 409.28 274.18 410 ;
    END
  END waddr_a_i[3]
  PIN waddr_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  275.42 409.28 275.62 410 ;
    END
  END waddr_a_i[4]
  PIN wdata_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  176.06 409.28 176.26 410 ;
    END
  END wdata_a_i[0]
  PIN wdata_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  276.86 409.28 277.06 410 ;
    END
  END wdata_a_i[10]
  PIN wdata_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  240.86 409.28 241.06 410 ;
    END
  END wdata_a_i[11]
  PIN wdata_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  223.58 409.28 223.78 410 ;
    END
  END wdata_a_i[12]
  PIN wdata_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  145.82 409.28 146.02 410 ;
    END
  END wdata_a_i[13]
  PIN wdata_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  201.98 409.28 202.18 410 ;
    END
  END wdata_a_i[14]
  PIN wdata_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  279.74 409.28 279.94 410 ;
    END
  END wdata_a_i[15]
  PIN wdata_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  281.18 409.28 281.38 410 ;
    END
  END wdata_a_i[16]
  PIN wdata_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  173.18 409.28 173.38 410 ;
    END
  END wdata_a_i[17]
  PIN wdata_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  258.14 409.28 258.34 410 ;
    END
  END wdata_a_i[18]
  PIN wdata_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  271.1 409.28 271.3 410 ;
    END
  END wdata_a_i[19]
  PIN wdata_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  163.1 409.28 163.3 410 ;
    END
  END wdata_a_i[1]
  PIN wdata_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  132.86 409.28 133.06 410 ;
    END
  END wdata_a_i[20]
  PIN wdata_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  249.5 409.28 249.7 410 ;
    END
  END wdata_a_i[21]
  PIN wdata_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  259.58 409.28 259.78 410 ;
    END
  END wdata_a_i[22]
  PIN wdata_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  282.62 409.28 282.82 410 ;
    END
  END wdata_a_i[23]
  PIN wdata_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  170.3 409.28 170.5 410 ;
    END
  END wdata_a_i[24]
  PIN wdata_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  144.38 409.28 144.58 410 ;
    END
  END wdata_a_i[25]
  PIN wdata_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  278.3 409.28 278.5 410 ;
    END
  END wdata_a_i[26]
  PIN wdata_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  284.06 409.28 284.26 410 ;
    END
  END wdata_a_i[27]
  PIN wdata_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  168.86 409.28 169.06 410 ;
    END
  END wdata_a_i[28]
  PIN wdata_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  250.94 409.28 251.14 410 ;
    END
  END wdata_a_i[29]
  PIN wdata_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  268.22 409.28 268.42 410 ;
    END
  END wdata_a_i[2]
  PIN wdata_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  158.78 409.28 158.98 410 ;
    END
  END wdata_a_i[30]
  PIN wdata_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  167.42 409.28 167.62 410 ;
    END
  END wdata_a_i[31]
  PIN wdata_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  272.54 409.28 272.74 410 ;
    END
  END wdata_a_i[3]
  PIN wdata_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  142.94 409.28 143.14 410 ;
    END
  END wdata_a_i[4]
  PIN wdata_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  194.78 409.28 194.98 410 ;
    END
  END wdata_a_i[5]
  PIN wdata_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  165.98 409.28 166.18 410 ;
    END
  END wdata_a_i[6]
  PIN wdata_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  261.02 409.28 261.22 410 ;
    END
  END wdata_a_i[7]
  PIN wdata_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  252.38 409.28 252.58 410 ;
    END
  END wdata_a_i[8]
  PIN wdata_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  285.5 409.28 285.7 410 ;
    END
  END wdata_a_i[9]
  PIN we_a_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  164.54 409.28 164.74 410 ;
    END
  END we_a_i
  OBS
    LAYER Metal1 ;
     RECT  5.28 7.34 404.64 404.68 ;
    LAYER Metal2 ;
     RECT  5.66 231.32 6.14 231.52 ;
     RECT  5.66 259.04 6.14 259.24 ;
     RECT  5.66 159.92 6.56 160.12 ;
     RECT  6.14 223.76 6.56 231.52 ;
     RECT  5.66 246.44 6.56 246.64 ;
     RECT  6.14 255.68 6.56 259.24 ;
     RECT  6.14 292.64 6.56 293.26 ;
     RECT  5.66 304.82 6.56 305.02 ;
     RECT  6.14 190.58 7.04 197.92 ;
     RECT  6.14 210.32 7.04 210.52 ;
     RECT  6.56 223.76 7.04 259.24 ;
     RECT  6.14 337.16 7.04 345.76 ;
     RECT  6.56 159.92 7.1 161.13 ;
     RECT  6.56 292.64 7.1 305.02 ;
     RECT  6.62 138.08 7.52 140.8 ;
     RECT  7.04 221.205 7.58 259.24 ;
     RECT  7.1 277.94 7.58 305.02 ;
     RECT  7.04 190.58 8 198.93 ;
     RECT  7.1 159.92 8.06 169.36 ;
     RECT  7.04 209.31 8.06 210.52 ;
     RECT  7.58 221.205 8.06 305.02 ;
     RECT  7.04 330.27 8.06 345.76 ;
     RECT  7.52 138.045 8.54 140.8 ;
     RECT  8.06 159.92 8.54 175.24 ;
     RECT  8 186.63 8.54 198.93 ;
     RECT  8.06 209.31 8.54 305.02 ;
     RECT  8.06 327.5 8.54 349.54 ;
     RECT  8.54 135.14 9.02 140.8 ;
     RECT  9.02 131.36 9.5 140.8 ;
     RECT  8.54 149.84 9.5 198.93 ;
     RECT  9.5 131.36 9.98 198.93 ;
     RECT  8.54 209.31 9.98 349.54 ;
     RECT  10.94 122.54 11.42 122.74 ;
     RECT  9.98 131.36 11.42 349.54 ;
     RECT  11.42 122.54 17.66 349.54 ;
     RECT  17.18 107 18.08 107.2 ;
     RECT  18.62 96.92 19.52 97.12 ;
     RECT  18.08 107 19.58 108.21 ;
     RECT  17.66 122.54 19.58 353.74 ;
     RECT  19.58 107 20.06 112.24 ;
     RECT  19.58 122.54 20.06 354.58 ;
     RECT  19.52 95.91 20.54 97.12 ;
     RECT  20.06 107 20.54 354.58 ;
     RECT  20.54 95.91 21.02 354.58 ;
     RECT  21.02 95.91 21.5 357.52 ;
     RECT  21.5 95.91 22.94 372.22 ;
     RECT  22.94 88.94 27.74 372.22 ;
     RECT  27.74 84.74 33.5 372.22 ;
     RECT  33.5 81.8 34.88 372.22 ;
     RECT  34.88 80.79 42.325 372.22 ;
     RECT  42.325 80.96 43.78 372.22 ;
     RECT  43.78 82.22 45.7 372.22 ;
     RECT  45.7 83.48 49.34 372.22 ;
     RECT  48.86 385.46 49.34 385.66 ;
     RECT  49.34 83.48 60.38 385.66 ;
     RECT  60.38 83.48 64.22 386.5 ;
     RECT  64.22 83.48 67.58 390.28 ;
     RECT  67.58 83.48 69.02 392.8 ;
     RECT  69.02 81.8 69.92 392.8 ;
     RECT  69.92 80.79 81.5 392.8 ;
     RECT  81.5 78.02 83.42 392.8 ;
     RECT  56.54 409.4 83.9 409.6 ;
     RECT  83.42 77.18 84.86 392.8 ;
     RECT  84.86 76.76 85.34 392.8 ;
     RECT  85.34 76.76 96.32 393.22 ;
     RECT  96.32 73.23 103.765 393.22 ;
     RECT  103.765 73.82 110.3 393.22 ;
     RECT  110.3 73.82 113.18 393.64 ;
     RECT  113.18 72.56 114.14 393.64 ;
     RECT  114.14 72.56 115.1 394.06 ;
     RECT  115.1 70.88 118.88 395.32 ;
     RECT  118.88 70.005 119.17 395.32 ;
     RECT  83.9 408.56 125.86 409.6 ;
     RECT  119.17 70.04 126.325 395.32 ;
     RECT  126.325 70.88 129.7 395.32 ;
     RECT  125.86 408.56 130.18 408.76 ;
     RECT  129.7 73.23 139.285 395.32 ;
     RECT  137.18 403.94 141.98 404.14 ;
     RECT  141.98 403.94 144.38 404.56 ;
     RECT  139.285 73.4 144.58 395.32 ;
     RECT  144.38 403.94 145.06 405.4 ;
     RECT  144.58 75.92 154.94 395.32 ;
     RECT  154.94 74.24 156.1 395.32 ;
     RECT  156.1 74.24 156.32 394.9 ;
     RECT  145.06 404.36 163.1 405.4 ;
     RECT  156.32 73.23 163.765 394.9 ;
     RECT  163.1 404.36 166.18 408.76 ;
     RECT  163.765 73.4 168.58 394.9 ;
     RECT  166.18 408.56 176.06 408.76 ;
     RECT  168.58 76.34 181.82 394.9 ;
     RECT  181.82 75.08 189.02 394.9 ;
     RECT  176.06 408.14 189.02 408.76 ;
     RECT  189.02 75.08 190.18 408.76 ;
     RECT  190.18 75.08 196.7 408.34 ;
     RECT  196.7 73.82 198.14 408.34 ;
     RECT  198.14 72.14 205.54 408.34 ;
     RECT  205.54 72.14 208.7 404.14 ;
     RECT  208.7 69.2 215.42 404.14 ;
     RECT  215.42 66.68 217.34 404.14 ;
     RECT  217.34 65.84 224.26 404.14 ;
     RECT  224.26 69.2 225.98 404.14 ;
     RECT  225.98 69.2 237.98 404.98 ;
     RECT  237.98 69.2 247.1 405.82 ;
     RECT  247.1 66.26 249.02 405.82 ;
     RECT  249.02 65.42 250.18 405.82 ;
     RECT  250.18 65.42 251.14 404.98 ;
     RECT  251.14 65.42 253.54 399.1 ;
     RECT  253.54 65.84 265.06 399.1 ;
     RECT  265.06 65.84 266.5 397.84 ;
     RECT  266.5 66.26 275.42 397.84 ;
     RECT  275.42 65 280.9 397.84 ;
     RECT  280.9 65 295.1 395.74 ;
     RECT  295.1 62.06 297.02 395.74 ;
     RECT  297.02 61.64 303.94 395.74 ;
     RECT  303.94 61.64 306.82 395.32 ;
     RECT  306.82 62.06 308.74 395.32 ;
     RECT  308.74 62.48 309.7 395.32 ;
     RECT  309.7 65.67 319.765 395.32 ;
     RECT  319.765 67.1 323.14 395.32 ;
     RECT  323.14 69.62 328.9 395.32 ;
     RECT  328.9 70.04 329.38 395.32 ;
     RECT  329.38 70.04 339.2 394.9 ;
     RECT  339.2 70.005 339.74 394.9 ;
     RECT  339.74 68.78 344.54 394.9 ;
     RECT  344.54 67.1 352.11 394.9 ;
     RECT  352.11 66.26 353.18 394.9 ;
     RECT  353.18 65.42 360.38 394.9 ;
     RECT  360.38 65 363.46 394.9 ;
     RECT  363.46 65 364.42 393.22 ;
     RECT  364.42 66.26 368.74 393.22 ;
     RECT  368.74 393.02 370.18 393.22 ;
     RECT  368.74 66.26 372.1 378.1 ;
     RECT  372.1 69.2 384.1 378.1 ;
     RECT  384.1 69.2 385.54 377.26 ;
     RECT  385.54 69.2 386.5 376 ;
     RECT  386.5 69.2 387.46 372.64 ;
     RECT  387.46 73.82 388.065 372.64 ;
     RECT  388.065 77.6 391.285 372.64 ;
     RECT  391.285 78.44 393.22 372.64 ;
     RECT  393.22 78.44 394.66 82.42 ;
     RECT  393.22 91.46 396.58 372.64 ;
     RECT  396.58 99.85 397.06 372.64 ;
     RECT  397.06 99.85 398.885 372.22 ;
     RECT  394.66 82.22 399.46 82.42 ;
     RECT  398.885 99.86 399.925 372.22 ;
     RECT  399.925 251.48 400.405 372.22 ;
     RECT  399.925 99.86 400.885 242.86 ;
     RECT  400.405 251.48 400.885 295.78 ;
     RECT  400.405 304.4 400.885 372.22 ;
     RECT  400.885 165.38 401.025 242.86 ;
     RECT  400.885 99.86 401.86 107.2 ;
     RECT  400.885 116.24 401.86 154.24 ;
     RECT  400.885 252.32 401.86 295.78 ;
     RECT  400.885 305.24 402.34 372.22 ;
     RECT  401.025 184.28 403.3 242.86 ;
     RECT  402.34 369.5 403.3 372.22 ;
     RECT  401.86 127.58 403.78 154.24 ;
     RECT  403.3 206.96 403.78 241.18 ;
     RECT  401.86 293.9 403.78 295.78 ;
     RECT  401.86 104.9 404.26 105.1 ;
     RECT  401.86 116.24 404.26 118.12 ;
     RECT  403.78 127.58 404.26 129.46 ;
     RECT  403.78 145.22 404.26 154.24 ;
     RECT  401.025 165.38 404.26 174.82 ;
     RECT  403.3 184.28 404.26 193.72 ;
     RECT  403.78 206.96 404.26 212.62 ;
     RECT  403.78 225.86 404.26 241.18 ;
     RECT  401.86 252.32 404.26 263.86 ;
     RECT  401.86 275 404.26 284.44 ;
     RECT  402.34 305.24 404.26 354.58 ;
    LAYER Metal3 ;
     RECT  299.42 61.64 299.62 62.06 ;
     RECT  299.42 62.06 308.74 62.48 ;
     RECT  296.06 62.48 309.7 64.7 ;
     RECT  295.58 64.7 309.7 65 ;
     RECT  280.7 65 309.7 65.42 ;
     RECT  360.38 65 360.58 65.42 ;
     RECT  275.9 65.42 309.7 65.84 ;
     RECT  358.46 65.42 361.54 65.84 ;
     RECT  224.06 65.84 224.26 66.26 ;
     RECT  249.02 65.42 253.54 66.26 ;
     RECT  275.9 65.84 312.58 66.26 ;
     RECT  355.1 65.84 361.54 66.26 ;
     RECT  219.74 66.26 224.26 66.68 ;
     RECT  275.9 66.26 313.06 66.68 ;
     RECT  273.5 66.68 316.42 67.1 ;
     RECT  352.7 66.26 361.54 67.1 ;
     RECT  344.54 67.1 361.54 68.78 ;
     RECT  218.3 66.68 224.26 69.2 ;
     RECT  246.14 66.26 253.54 69.2 ;
     RECT  218.3 69.2 253.54 69.62 ;
     RECT  273.02 67.1 320.74 69.62 ;
     RECT  371.9 66.26 372.1 69.62 ;
     RECT  387.26 69.2 387.46 69.62 ;
     RECT  119.9 69.62 120.1 70.04 ;
     RECT  218.3 69.62 263.14 70.04 ;
     RECT  273.02 69.62 328.9 70.04 ;
     RECT  339.74 68.78 361.54 70.04 ;
     RECT  217.82 70.04 263.14 70.88 ;
     RECT  117.98 70.04 126.34 72.98 ;
     RECT  113.18 72.98 126.34 73.4 ;
     RECT  214.94 70.88 263.14 73.4 ;
     RECT  273.02 70.04 361.54 73.4 ;
     RECT  371.9 69.62 387.46 73.4 ;
     RECT  96.38 73.4 96.58 73.82 ;
     RECT  113.18 73.4 129.7 73.82 ;
     RECT  144.38 73.4 144.58 73.82 ;
     RECT  168.38 73.4 168.58 73.82 ;
     RECT  209.18 73.4 387.46 73.82 ;
     RECT  96.38 73.82 144.58 74.24 ;
     RECT  198.14 72.14 198.34 74.24 ;
     RECT  162.14 73.82 168.58 74.66 ;
     RECT  198.14 74.24 198.82 74.66 ;
     RECT  209.18 73.82 387.94 74.66 ;
     RECT  95.42 74.24 144.58 75.92 ;
     RECT  161.18 74.66 168.58 75.92 ;
     RECT  181.82 75.08 182.02 76.34 ;
     RECT  198.14 74.66 387.94 76.34 ;
     RECT  95.42 75.92 168.58 76.76 ;
     RECT  91.58 76.76 168.58 77.18 ;
     RECT  181.82 76.34 387.94 77.18 ;
     RECT  83.42 77.18 387.94 78.02 ;
     RECT  81.5 78.02 387.94 78.44 ;
     RECT  81.5 78.44 388.9 80.96 ;
     RECT  43.58 80.96 43.78 81.38 ;
     RECT  77.66 80.96 388.9 81.38 ;
     RECT  37.34 81.38 43.78 81.8 ;
     RECT  70.94 81.38 388.9 83.9 ;
     RECT  33.5 81.8 43.78 84.32 ;
     RECT  33.02 84.32 43.78 84.74 ;
     RECT  67.58 83.9 388.9 85.16 ;
     RECT  399.26 82.22 399.46 85.16 ;
     RECT  27.74 84.74 52.9 86 ;
     RECT  66.14 85.16 399.46 86 ;
     RECT  27.74 86 399.46 88.94 ;
     RECT  22.94 88.94 399.46 96.5 ;
     RECT  20.54 96.5 399.46 99.64 ;
     RECT  21.5 99.64 399.46 99.86 ;
     RECT  21.5 99.86 401.86 114.56 ;
     RECT  20.06 114.56 401.86 122.12 ;
     RECT  12.86 122.12 401.86 122.54 ;
     RECT  11.42 122.54 401.86 124.84 ;
     RECT  11.42 124.84 398.02 134.5 ;
     RECT  11.42 134.5 396.1 135.14 ;
     RECT  8.54 135.14 396.1 137.44 ;
     RECT  8.54 137.44 395.62 137.86 ;
     RECT  9.98 137.86 395.62 149.42 ;
     RECT  8.06 149.42 395.62 153.2 ;
     RECT  8.06 153.2 397.54 161.6 ;
     RECT  8.06 161.6 404.26 169.16 ;
     RECT  7.1 169.16 404.26 172.3 ;
     RECT  7.1 172.3 403.3 174.82 ;
     RECT  7.1 174.82 401.38 187 ;
     RECT  7.58 187 401.38 190.78 ;
     RECT  7.58 190.78 399.94 192.46 ;
     RECT  7.58 192.46 399.46 194.98 ;
     RECT  8.06 194.98 399.46 201.7 ;
     RECT  8.06 201.7 398.98 205.06 ;
     RECT  8.06 205.06 398.02 211.78 ;
     RECT  8.06 211.78 397.54 221.24 ;
     RECT  6.14 221.24 397.54 228.8 ;
     RECT  5.66 228.8 397.54 251.9 ;
     RECT  5.66 251.9 398.02 252.32 ;
     RECT  5.66 252.32 401.38 258.82 ;
     RECT  5.66 258.82 398.02 259.24 ;
     RECT  7.1 259.24 398.02 280.88 ;
     RECT  7.1 280.88 400.9 296.84 ;
     RECT  5.66 296.84 400.9 299.56 ;
     RECT  5.66 299.56 399.46 300.82 ;
     RECT  5.66 300.82 398.5 305.02 ;
     RECT  10.46 305.02 398.5 315.74 ;
     RECT  8.54 315.74 398.5 316.58 ;
     RECT  8.54 316.58 398.98 319.52 ;
     RECT  8.06 319.52 398.98 320.36 ;
     RECT  8.06 320.36 404.26 330.86 ;
     RECT  6.14 330.86 404.26 334.42 ;
     RECT  6.14 334.42 400.42 345.76 ;
     RECT  7.58 345.76 400.42 346.18 ;
     RECT  9.5 346.18 400.42 348.92 ;
     RECT  9.5 348.92 401.38 349.12 ;
     RECT  11.42 349.12 401.38 350.38 ;
     RECT  19.58 350.38 401.38 353.74 ;
     RECT  21.5 353.74 401.38 360.46 ;
     RECT  21.5 360.46 400.42 362.56 ;
     RECT  21.5 362.56 397.06 368.44 ;
     RECT  21.5 368.44 26.5 369.28 ;
     RECT  43.1 368.44 397.06 369.28 ;
     RECT  46.46 369.28 397.06 370.54 ;
     RECT  48.86 370.54 397.06 371.8 ;
     RECT  21.5 369.28 21.7 372.22 ;
     RECT  81.98 371.8 397.06 372.64 ;
     RECT  48.86 371.8 72.1 373.06 ;
     RECT  81.98 372.64 388.42 373.06 ;
     RECT  104.06 373.06 386.98 373.48 ;
     RECT  83.9 373.06 89.38 373.9 ;
     RECT  110.3 373.48 386.98 375.16 ;
     RECT  110.3 375.16 386.5 376 ;
     RECT  110.3 376 384.58 376.42 ;
     RECT  383.42 376.42 384.1 377.26 ;
     RECT  383.9 377.26 384.1 378.1 ;
     RECT  110.3 376.42 370.18 379.78 ;
     RECT  351.74 379.78 370.18 380.2 ;
     RECT  110.3 379.78 338.98 382.72 ;
     RECT  321.98 382.72 338.98 383.14 ;
     RECT  110.3 382.72 311.62 383.56 ;
     RECT  48.86 373.06 67.78 385.66 ;
     RECT  322.94 383.14 338.98 386.08 ;
     RECT  110.3 383.56 311.14 386.92 ;
     RECT  322.94 386.08 334.18 388.6 ;
     RECT  56.54 385.66 67.78 390.28 ;
     RECT  124.22 386.92 311.14 390.28 ;
     RECT  124.22 390.28 303.94 392.38 ;
     RECT  67.58 390.28 67.78 392.8 ;
     RECT  83.9 373.9 85.54 393.22 ;
     RECT  354.14 380.2 370.18 393.22 ;
     RECT  110.3 386.92 114.34 393.64 ;
     RECT  322.94 388.6 329.38 393.64 ;
     RECT  114.14 393.64 114.34 394.06 ;
     RECT  326.78 393.64 329.38 394.06 ;
     RECT  354.14 393.22 363.46 394.48 ;
     RECT  363.26 394.48 363.46 394.9 ;
     RECT  329.18 394.06 329.38 395.32 ;
     RECT  303.74 392.38 303.94 395.74 ;
     RECT  83.9 393.22 84.1 408.76 ;
     RECT  124.22 392.38 287.14 409.5 ;
     RECT  56.54 390.28 56.74 409.6 ;
     RECT  131.9 409.5 135.46 409.6 ;
     RECT  156.38 409.5 157.06 409.6 ;
     RECT  173.66 409.5 185.86 409.6 ;
     RECT  203.9 409.5 217.54 409.6 ;
     RECT  232.7 409.5 233.38 409.6 ;
     RECT  248.54 409.5 270.82 409.6 ;
     RECT  283.1 409.5 285.22 409.6 ;
    LAYER Metal4 ;
     RECT  14.3 300.62 15.26 300.82 ;
     RECT  9.5 258.62 16.22 258.82 ;
     RECT  9.98 285.5 16.22 285.7 ;
     RECT  14.78 201.92 17.86 202.12 ;
     RECT  17.66 315.74 19.58 315.94 ;
     RECT  19.58 315.74 20.06 323.5 ;
     RECT  13.34 126.74 21.7 126.94 ;
     RECT  15.26 300.2 21.98 300.82 ;
     RECT  20.06 315.74 22.66 323.92 ;
     RECT  15.26 233 22.94 233.2 ;
     RECT  21.98 342.2 23.42 342.4 ;
     RECT  16.22 258.62 23.62 263.02 ;
     RECT  23.42 342.2 25.82 349.96 ;
     RECT  19.1 243.92 26.78 244.12 ;
     RECT  22.94 232.58 27.74 233.2 ;
     RECT  25.82 334.22 27.94 349.96 ;
     RECT  21.98 300.2 28.7 304.18 ;
     RECT  22.66 318.26 28.7 323.92 ;
     RECT  27.94 334.22 28.7 346.6 ;
     RECT  16.22 281.3 28.9 285.7 ;
     RECT  27.74 228.8 31.78 233.2 ;
     RECT  28.9 285.5 33.02 285.7 ;
     RECT  28.7 296.42 33.02 304.18 ;
     RECT  33.02 285.5 33.5 304.18 ;
     RECT  33.5 285.5 33.98 308.8 ;
     RECT  28.7 318.26 33.98 346.6 ;
     RECT  33.02 104.06 34.46 104.26 ;
     RECT  33.98 285.5 34.66 346.6 ;
     RECT  27.26 145.22 34.94 145.42 ;
     RECT  34.94 141.44 35.42 145.42 ;
     RECT  33.02 269.54 35.42 269.74 ;
     RECT  32.06 213.26 36.38 213.46 ;
     RECT  34.94 122.12 37.34 122.32 ;
     RECT  35.42 141.44 37.82 153.4 ;
     RECT  26.78 243.92 37.82 253.78 ;
     RECT  35.42 265.34 37.82 269.74 ;
     RECT  37.82 141.44 38.78 157.18 ;
     RECT  36.38 205.7 38.78 213.46 ;
     RECT  37.82 243.92 38.98 269.74 ;
     RECT  34.66 285.5 38.98 330.22 ;
     RECT  31.78 228.8 39.46 232.78 ;
     RECT  38.98 259.88 39.74 269.74 ;
     RECT  38.98 243.92 39.94 251.26 ;
     RECT  34.66 338.84 40.22 346.6 ;
     RECT  38.98 285.5 40.42 328.12 ;
     RECT  39.74 259.88 40.7 274.36 ;
     RECT  40.42 285.5 40.7 308.8 ;
     RECT  38.78 204.86 41.38 213.46 ;
     RECT  39.94 247.28 41.38 251.26 ;
     RECT  40.7 259.88 41.38 308.8 ;
     RECT  40.22 338.84 41.38 352.48 ;
     RECT  37.34 122.12 41.66 123.16 ;
     RECT  34.46 99.86 42.34 104.26 ;
     RECT  41.38 259.88 42.34 302.5 ;
     RECT  40.42 318.26 42.82 328.12 ;
     RECT  41.66 115.4 43.1 123.16 ;
     RECT  42.82 318.26 43.3 327.28 ;
     RECT  42.34 262.82 43.78 269.74 ;
     RECT  43.3 318.26 43.78 323.5 ;
     RECT  43.1 115.4 44.26 126.94 ;
     RECT  38.78 138.92 44.26 157.18 ;
     RECT  42.34 281.72 44.26 302.5 ;
     RECT  41.38 209.48 44.54 213.46 ;
     RECT  39.46 232.58 44.74 232.78 ;
     RECT  44.26 115.4 45.22 116.02 ;
     RECT  43.78 318.26 45.22 323.08 ;
     RECT  44.54 209.48 45.7 216.82 ;
     RECT  44.26 281.72 46.18 281.92 ;
     RECT  42.34 99.86 47.14 100.06 ;
     RECT  44.26 126.74 47.14 126.94 ;
     RECT  41.66 171.68 47.14 171.88 ;
     RECT  44.26 141.44 47.62 157.18 ;
     RECT  41.38 341.78 47.62 352.48 ;
     RECT  45.7 209.48 49.06 209.68 ;
     RECT  45.22 115.4 49.54 115.6 ;
     RECT  47.62 352.28 50.02 352.48 ;
     RECT  41.38 251.06 50.3 251.26 ;
     RECT  44.26 292.64 50.3 302.5 ;
     RECT  48.38 165.8 50.5 166 ;
     RECT  50.3 242.66 50.5 251.26 ;
     RECT  43.78 262.82 50.5 265.54 ;
     RECT  50.5 242.66 50.78 250.84 ;
     RECT  48.38 221.66 50.98 224.8 ;
     RECT  47.62 341.78 51.74 342.82 ;
     RECT  52.22 100.28 53.66 100.48 ;
     RECT  50.3 292.64 53.86 306.28 ;
     RECT  50.78 240.56 54.62 250.84 ;
     RECT  53.66 100.28 56.26 108.04 ;
     RECT  54.62 129.26 57.02 129.46 ;
     RECT  47.62 141.44 57.02 147.1 ;
     RECT  51.74 338.42 57.5 342.82 ;
     RECT  53.18 364.88 57.98 365.08 ;
     RECT  55.58 202.34 58.46 202.54 ;
     RECT  50.98 221.66 58.94 221.86 ;
     RECT  58.94 221.24 59.14 221.86 ;
     RECT  54.62 284.66 60.38 284.86 ;
     RECT  57.5 338.42 60.38 344.5 ;
     RECT  57.98 268.7 60.86 268.9 ;
     RECT  57.02 129.26 61.06 147.1 ;
     RECT  60.38 280.88 62.02 284.86 ;
     RECT  57.98 364.46 62.3 365.08 ;
     RECT  54.62 237.62 63.74 250.84 ;
     RECT  60.86 268.7 64.22 270.16 ;
     RECT  60.38 338.42 64.22 349.96 ;
     RECT  62.3 364.46 64.42 370.54 ;
     RECT  53.86 296.42 64.7 306.28 ;
     RECT  62.02 280.88 64.9 281.08 ;
     RECT  64.7 296.42 65.18 310.9 ;
     RECT  45.22 322.88 65.18 323.08 ;
     RECT  65.18 296.42 68.26 323.08 ;
     RECT  63.74 237.62 69.02 255.04 ;
     RECT  69.02 232.58 69.22 255.04 ;
     RECT  65.66 160.76 69.98 160.96 ;
     RECT  56.26 101.12 70.94 104.26 ;
     RECT  64.42 364.46 71.14 365.08 ;
     RECT  69.98 160.76 72.58 165.16 ;
     RECT  64.22 266.18 73.34 270.16 ;
     RECT  72.86 281.72 73.34 281.92 ;
     RECT  68.54 175.88 73.54 176.08 ;
     RECT  61.06 130.94 73.82 147.1 ;
     RECT  58.46 198.56 74.3 202.54 ;
     RECT  64.22 334.64 74.5 349.96 ;
     RECT  74.3 198.56 74.78 202.96 ;
     RECT  74.78 198.56 75.26 205.9 ;
     RECT  74.5 348.5 75.26 349.96 ;
     RECT  69.22 232.58 76.42 250.84 ;
     RECT  68.26 296.42 76.42 319.3 ;
     RECT  71.9 221.24 76.9 221.44 ;
     RECT  70.94 100.28 77.66 104.26 ;
     RECT  74.5 334.64 77.86 338.62 ;
     RECT  63.26 121.7 79.1 121.9 ;
     RECT  73.82 130.52 79.1 147.1 ;
     RECT  79.1 121.7 79.3 147.1 ;
     RECT  77.66 99.86 80.06 104.26 ;
     RECT  76.42 298.94 80.26 319.3 ;
     RECT  75.26 194.78 80.74 205.9 ;
     RECT  76.42 232.58 81.7 232.78 ;
     RECT  71.14 364.46 81.7 364.66 ;
     RECT  73.34 266.18 81.98 281.92 ;
     RECT  81.98 168.32 82.46 168.52 ;
     RECT  80.74 198.56 82.66 205.9 ;
     RECT  76.42 242.66 82.66 250.84 ;
     RECT  80.26 319.1 82.94 319.3 ;
     RECT  81.98 262.82 83.42 281.92 ;
     RECT  82.66 243.08 83.62 250.84 ;
     RECT  82.46 164.54 85.06 168.52 ;
     RECT  77.86 338.42 85.06 338.62 ;
     RECT  83.42 259.88 86.02 281.92 ;
     RECT  86.02 266.18 87.46 281.92 ;
     RECT  79.3 136.82 88.9 147.1 ;
     RECT  75.26 348.5 89.66 353.74 ;
     RECT  82.94 319.1 90.14 319.72 ;
     RECT  90.14 319.1 90.34 326.86 ;
     RECT  82.66 198.56 90.82 202.54 ;
     RECT  79.3 121.7 91.3 123.16 ;
     RECT  88.9 137.24 91.3 147.1 ;
     RECT  80.06 99.86 92.06 104.68 ;
     RECT  85.06 168.32 92.06 168.52 ;
     RECT  92.06 99.86 92.26 107.2 ;
     RECT  83.62 243.08 92.26 247.48 ;
     RECT  80.26 298.94 92.26 307.96 ;
     RECT  89.66 348.5 92.26 357.52 ;
     RECT  92.26 307.76 93.02 307.96 ;
     RECT  91.3 137.66 93.22 147.1 ;
     RECT  92.06 168.32 93.22 170.2 ;
     RECT  87.46 266.18 93.22 277.72 ;
     RECT  92.26 357.32 93.7 357.52 ;
     RECT  93.22 137.66 94.18 142.06 ;
     RECT  93.02 197.72 94.94 197.92 ;
     RECT  85.34 216.2 94.94 216.4 ;
     RECT  90.34 326.66 95.14 326.86 ;
     RECT  93.02 307.76 96.1 314.26 ;
     RECT  94.94 209.9 96.58 216.4 ;
     RECT  91.3 122.96 98.98 123.16 ;
     RECT  94.18 141.86 99.46 142.06 ;
     RECT  90.14 288.86 99.74 289.06 ;
     RECT  93.22 266.18 99.94 266.38 ;
     RECT  93.22 168.32 100.42 168.52 ;
     RECT  93.22 277.52 100.7 277.72 ;
     RECT  99.74 288.86 100.7 289.48 ;
     RECT  92.26 298.94 100.7 299.14 ;
     RECT  100.7 277.52 100.9 299.14 ;
     RECT  92.26 348.5 100.9 348.7 ;
     RECT  96.58 216.2 102.34 216.4 ;
     RECT  92.26 104.06 103.3 107.2 ;
     RECT  92.26 243.08 103.58 246.64 ;
     RECT  101.66 268.7 103.78 268.9 ;
     RECT  103.58 242.24 104.06 246.64 ;
     RECT  104.06 242.24 105.22 259.24 ;
     RECT  94.94 195.62 105.5 197.92 ;
     RECT  104.06 92.3 105.98 92.5 ;
     RECT  102.14 164.54 107.42 168.1 ;
     RECT  107.42 163.28 107.62 168.1 ;
     RECT  105.22 242.24 107.62 250.42 ;
     RECT  105.5 111.62 107.9 111.82 ;
     RECT  106.46 130.52 108.38 130.72 ;
     RECT  105.5 195.62 108.38 202.12 ;
     RECT  108.38 190.58 110.98 202.12 ;
     RECT  105.98 91.46 112.7 92.5 ;
     RECT  107.62 164.54 112.7 168.1 ;
     RECT  112.7 164.54 112.9 176.08 ;
     RECT  112.7 91.46 113.18 100.48 ;
     RECT  107.9 111.62 113.18 115.18 ;
     RECT  108.38 130.52 113.38 134.5 ;
     RECT  100.9 285.08 115.1 297.46 ;
     RECT  110.78 322.88 115.1 323.08 ;
     RECT  107.62 242.24 115.78 242.86 ;
     RECT  113.18 91.46 117.22 115.18 ;
     RECT  117.02 217.46 117.5 217.66 ;
     RECT  111.74 228.8 117.5 229 ;
     RECT  110.98 201.92 118.66 202.12 ;
     RECT  115.1 315.74 118.94 323.08 ;
     RECT  115.1 285.08 120.1 300.4 ;
     RECT  117.5 217.46 120.58 229 ;
     RECT  118.94 315.74 120.58 325.6 ;
     RECT  118.94 341.36 120.58 346.18 ;
     RECT  113.38 130.52 121.54 130.72 ;
     RECT  120.58 228.8 121.54 229 ;
     RECT  112.9 168.32 122.5 176.08 ;
     RECT  122.5 168.32 123.94 172.3 ;
     RECT  117.98 273.74 124.22 273.94 ;
     RECT  120.1 288.44 124.22 300.4 ;
     RECT  120.58 315.74 124.22 323.08 ;
     RECT  120.58 341.36 125.38 345.34 ;
     RECT  117.22 99.86 125.86 115.18 ;
     RECT  121.34 360.68 126.14 360.88 ;
     RECT  123.94 168.32 127.78 168.52 ;
     RECT  110.98 190.58 129.02 190.78 ;
     RECT  119.42 247.7 129.02 247.9 ;
     RECT  105.22 259.04 129.02 259.24 ;
     RECT  129.02 247.7 129.22 259.24 ;
     RECT  125.86 99.86 130.18 111.82 ;
     RECT  124.22 288.44 130.18 323.08 ;
     RECT  124.22 134.3 130.94 134.5 ;
     RECT  127.58 236.78 131.62 236.98 ;
     RECT  130.18 100.28 132.1 111.82 ;
     RECT  130.94 126.74 132.86 134.5 ;
     RECT  123.26 73.82 133.06 74.02 ;
     RECT  130.18 288.44 133.54 313.42 ;
     RECT  126.14 356.48 133.54 360.88 ;
     RECT  125.38 341.36 133.82 341.56 ;
     RECT  133.54 356.48 133.82 357.52 ;
     RECT  124.22 273.74 134.3 277.72 ;
     RECT  133.54 288.44 134.3 300.82 ;
     RECT  132.86 126.74 135.26 138.7 ;
     RECT  127.58 156.56 135.74 156.76 ;
     RECT  130.18 322.88 135.74 323.08 ;
     RECT  133.82 341.36 136.42 357.52 ;
     RECT  132.1 100.28 136.9 104.26 ;
     RECT  129.02 190.58 137.18 199.18 ;
     RECT  136.9 100.28 137.86 103.84 ;
     RECT  120.58 217.46 137.86 217.66 ;
     RECT  137.18 190.58 138.34 207.16 ;
     RECT  134.3 273.74 138.82 300.82 ;
     RECT  135.74 322.88 138.82 323.5 ;
     RECT  138.82 273.74 140.26 273.94 ;
     RECT  129.22 247.7 140.74 252.52 ;
     RECT  129.02 375.8 141.02 376 ;
     RECT  136.42 341.36 142.94 341.98 ;
     RECT  140.74 247.7 143.14 247.9 ;
     RECT  138.34 190.58 143.62 202.54 ;
     RECT  142.94 338 143.62 341.98 ;
     RECT  135.74 149.42 144.1 156.76 ;
     RECT  135.26 118.76 144.38 138.7 ;
     RECT  143.42 245.18 144.38 247.48 ;
     RECT  143.62 338 144.86 338.2 ;
     RECT  144.38 114.56 146.02 138.7 ;
     RECT  144.1 156.56 146.02 156.76 ;
     RECT  144.38 240.98 146.02 247.48 ;
     RECT  145.34 272.9 146.78 273.1 ;
     RECT  139.1 88.52 147.46 88.72 ;
     RECT  137.86 100.28 147.94 100.48 ;
     RECT  142.46 174.62 148.22 174.82 ;
     RECT  146.02 114.56 148.9 134.5 ;
     RECT  138.82 323.3 148.9 323.5 ;
     RECT  148.22 174.62 149.38 179.02 ;
     RECT  148.9 134.3 149.86 134.5 ;
     RECT  141.02 368.24 149.86 376 ;
     RECT  143.62 198.14 150.34 202.54 ;
     RECT  150.34 201.08 150.82 202.54 ;
     RECT  146.78 266.6 151.1 273.1 ;
     RECT  138.82 285.92 151.1 300.82 ;
     RECT  133.54 310.7 151.1 313.42 ;
     RECT  148.9 114.56 151.3 123.16 ;
     RECT  150.82 201.08 151.3 201.7 ;
     RECT  136.42 352.28 151.58 352.48 ;
     RECT  146.02 245.18 152.06 247.48 ;
     RECT  152.06 245.18 152.54 251.68 ;
     RECT  151.1 265.76 152.54 313.42 ;
     RECT  144.86 334.64 153.02 338.2 ;
     RECT  151.58 352.28 153.02 358.78 ;
     RECT  153.02 334.64 153.7 358.78 ;
     RECT  149.86 375.8 153.7 376 ;
     RECT  152.54 245.18 154.18 313.42 ;
     RECT  153.7 337.58 154.46 358.78 ;
     RECT  154.18 270.38 155.42 313.42 ;
     RECT  155.42 270.38 155.62 319.72 ;
     RECT  154.46 337.58 156.1 359.2 ;
     RECT  154.18 245.18 156.38 259.24 ;
     RECT  152.06 103.64 157.34 103.84 ;
     RECT  156.38 240.98 157.54 259.24 ;
     RECT  157.54 245.18 158.02 259.24 ;
     RECT  155.62 281.3 158.02 319.72 ;
     RECT  157.34 99.44 158.5 103.84 ;
     RECT  151.1 210.32 158.98 210.52 ;
     RECT  153.98 84.74 159.94 84.94 ;
     RECT  155.42 191 161.18 191.2 ;
     RECT  151.3 201.08 161.18 201.28 ;
     RECT  158.02 283.4 162.62 319.72 ;
     RECT  159.26 217.04 163.1 217.24 ;
     RECT  161.18 88.94 163.78 89.14 ;
     RECT  163.1 138.08 164.06 138.28 ;
     RECT  161.18 191 164.06 201.28 ;
     RECT  151.3 122.96 164.74 123.16 ;
     RECT  152.54 149.42 165.02 149.62 ;
     RECT  160.7 390.92 165.02 391.12 ;
     RECT  163.1 217.04 165.22 222.28 ;
     RECT  164.06 189.32 167.14 201.28 ;
     RECT  165.02 149.42 167.62 153.82 ;
     RECT  155.62 270.38 168.86 270.58 ;
     RECT  168.86 270.38 169.34 273.52 ;
     RECT  156.1 338 169.34 357.52 ;
     RECT  158.5 99.44 170.78 100.06 ;
     RECT  158.02 245.6 171.74 259.24 ;
     RECT  169.34 269.12 171.74 273.52 ;
     RECT  163.58 173.36 172.22 173.56 ;
     RECT  167.14 189.32 172.22 198.34 ;
     RECT  172.22 173.36 172.42 198.34 ;
     RECT  165.02 390.92 173.18 393.64 ;
     RECT  171.74 245.6 174.14 273.52 ;
     RECT  162.62 283.4 174.14 323.5 ;
     RECT  165.22 217.04 174.82 219.76 ;
     RECT  164.06 136.4 175.1 138.28 ;
     RECT  175.1 130.1 175.3 138.28 ;
     RECT  174.14 245.6 175.3 323.5 ;
     RECT  174.82 217.04 175.58 217.24 ;
     RECT  170.78 99.44 175.78 100.48 ;
     RECT  175.78 99.86 176.54 100.48 ;
     RECT  175.58 210.32 176.54 217.24 ;
     RECT  176.54 99.86 176.74 100.9 ;
     RECT  167.62 153.62 176.74 153.82 ;
     RECT  175.3 272.9 176.74 323.5 ;
     RECT  168.38 77.6 177.22 77.8 ;
     RECT  165.5 368.24 177.7 368.44 ;
     RECT  176.74 99.86 179.14 100.06 ;
     RECT  172.42 181.34 179.9 198.34 ;
     RECT  176.54 209.9 179.9 217.24 ;
     RECT  179.9 181.34 181.06 217.24 ;
     RECT  169.34 337.16 182.98 357.52 ;
     RECT  175.3 245.6 183.94 263.44 ;
     RECT  183.74 408.98 183.94 409.6 ;
     RECT  181.06 181.34 185.38 195.4 ;
     RECT  176.74 277.1 186.14 323.5 ;
     RECT  178.46 231.74 186.82 231.94 ;
     RECT  183.94 263.24 186.82 263.44 ;
     RECT  181.06 209.9 187.58 217.24 ;
     RECT  186.14 145.64 187.78 145.84 ;
     RECT  187.58 209.9 187.78 224.8 ;
     RECT  186.14 272.9 187.78 323.5 ;
     RECT  183.94 245.6 188.54 251.26 ;
     RECT  175.1 164.12 189.5 164.32 ;
     RECT  188.54 240.98 190.18 251.26 ;
     RECT  187.78 209.9 190.66 213.46 ;
     RECT  182.98 337.16 190.66 337.36 ;
     RECT  190.66 209.9 191.14 210.52 ;
     RECT  187.78 301.04 191.14 323.5 ;
     RECT  175.3 130.1 191.62 130.3 ;
     RECT  187.78 224.6 192.1 224.8 ;
     RECT  191.14 301.04 192.1 315.94 ;
     RECT  182.98 345.98 192.58 353.74 ;
     RECT  189.5 156.56 193.06 164.32 ;
     RECT  192.58 345.98 193.06 346.18 ;
     RECT  190.18 245.6 193.54 251.26 ;
     RECT  186.14 98.6 194.02 98.8 ;
     RECT  187.78 272.9 194.3 289.48 ;
     RECT  193.06 164.12 194.5 164.32 ;
     RECT  194.3 269.96 195.26 289.48 ;
     RECT  191.14 209.9 195.94 210.1 ;
     RECT  193.54 247.7 196.42 251.26 ;
     RECT  190.94 84.74 197.86 84.94 ;
     RECT  196.42 248.12 198.34 251.26 ;
     RECT  195.26 130.94 198.82 131.14 ;
     RECT  192.1 301.04 198.82 305.86 ;
     RECT  185.38 181.34 199.3 191.62 ;
     RECT  196.22 149.84 199.78 150.04 ;
     RECT  192.1 315.74 199.78 315.94 ;
     RECT  198.82 301.04 201.22 302.08 ;
     RECT  199.3 181.34 201.7 189.52 ;
     RECT  198.34 251.06 201.7 251.26 ;
     RECT  195.26 269.54 201.7 289.48 ;
     RECT  201.7 275 203.9 289.48 ;
     RECT  203.9 275 205.06 293.68 ;
     RECT  203.9 353.12 205.34 357.52 ;
     RECT  201.5 338 205.54 338.2 ;
     RECT  201.5 217.04 206.02 217.24 ;
     RECT  204.38 251.48 206.02 252.1 ;
     RECT  202.46 225.86 206.78 226.06 ;
     RECT  206.78 225.86 207.26 228.16 ;
     RECT  205.06 275 207.46 288.64 ;
     RECT  206.78 252.74 209.66 258.82 ;
     RECT  209.66 252.74 210.14 264.7 ;
     RECT  202.46 123.38 212.74 123.58 ;
     RECT  209.18 194.36 213.98 194.56 ;
     RECT  207.26 217.46 214.46 228.16 ;
     RECT  214.46 214.52 214.94 228.16 ;
     RECT  213.98 194.36 215.42 200.86 ;
     RECT  214.94 214.1 215.42 228.16 ;
     RECT  202.94 318.68 215.42 318.88 ;
     RECT  215.42 194.36 215.62 228.16 ;
     RECT  210.14 252.74 215.62 266.8 ;
     RECT  205.34 352.28 215.62 357.52 ;
     RECT  215.42 318.68 215.9 326.02 ;
     RECT  207.46 283.4 216.38 288.64 ;
     RECT  215.9 317.42 216.38 326.02 ;
     RECT  215.62 252.74 216.58 265.12 ;
     RECT  216.38 283.4 217.34 291.16 ;
     RECT  209.18 89.36 217.82 89.56 ;
     RECT  217.34 114.98 218.78 115.18 ;
     RECT  217.34 282.98 218.78 291.16 ;
     RECT  216.38 317.42 218.78 331.06 ;
     RECT  218.78 282.98 220.22 296.2 ;
     RECT  220.22 281.3 220.42 296.2 ;
     RECT  218.78 314.48 220.7 331.06 ;
     RECT  215.62 194.36 221.38 222.7 ;
     RECT  216.58 252.74 222.82 258.82 ;
     RECT  222.82 252.74 223.58 256.72 ;
     RECT  221.38 215.36 224.26 222.7 ;
     RECT  207.26 342.2 226.94 342.4 ;
     RECT  221.38 194.36 227.14 200.86 ;
     RECT  215.62 357.32 227.62 357.52 ;
     RECT  224.26 215.36 228.1 222.28 ;
     RECT  223.58 239.72 228.1 256.72 ;
     RECT  220.7 307.34 228.1 331.06 ;
     RECT  173.18 390.92 228.38 395.74 ;
     RECT  205.34 135.14 228.86 135.34 ;
     RECT  218.78 107.42 229.06 115.18 ;
     RECT  226.94 341.78 229.06 342.4 ;
     RECT  217.82 89.36 230.02 96.28 ;
     RECT  229.06 342.2 230.02 342.4 ;
     RECT  203.42 179.66 230.3 179.86 ;
     RECT  228.1 239.72 230.78 239.92 ;
     RECT  230.3 174.62 231.26 179.86 ;
     RECT  228.1 307.76 231.26 331.06 ;
     RECT  230.02 96.08 231.46 96.28 ;
     RECT  228.1 218.3 231.46 222.28 ;
     RECT  231.46 218.3 232.42 218.5 ;
     RECT  228.1 252.74 233.18 256.72 ;
     RECT  220.42 281.3 233.66 289.06 ;
     RECT  227.14 194.36 233.86 194.56 ;
     RECT  233.18 252.74 234.62 262.6 ;
     RECT  231.26 174.62 236.74 183.64 ;
     RECT  230.78 235.52 237.5 239.92 ;
     RECT  228.86 130.94 237.98 135.34 ;
     RECT  220.22 150.68 237.98 150.88 ;
     RECT  229.06 114.98 238.46 115.18 ;
     RECT  233.66 279.2 238.46 289.48 ;
     RECT  231.26 307.76 238.46 331.48 ;
     RECT  234.62 252.74 238.66 267.64 ;
     RECT  238.46 112.04 238.94 115.18 ;
     RECT  238.46 279.2 239.42 293.68 ;
     RECT  238.46 307.76 240.38 334.42 ;
     RECT  236.74 175.88 240.58 183.64 ;
     RECT  239.42 279.2 240.58 297.46 ;
     RECT  237.98 130.1 241.06 135.34 ;
     RECT  240.58 175.88 241.06 183.22 ;
     RECT  227.42 368.24 241.34 368.44 ;
     RECT  228.38 384.2 241.34 395.74 ;
     RECT  241.06 175.88 241.54 179.86 ;
     RECT  241.34 368.24 241.54 395.74 ;
     RECT  237.5 235.52 241.82 244.12 ;
     RECT  240.58 279.2 242.3 293.68 ;
     RECT  241.06 130.1 242.5 131.14 ;
     RECT  241.82 228.38 242.5 244.12 ;
     RECT  238.94 111.2 243.26 115.18 ;
     RECT  242.3 277.52 243.46 293.68 ;
     RECT  238.66 252.74 244.22 265.96 ;
     RECT  240.38 307.34 244.22 334.42 ;
     RECT  244.22 247.7 246.34 265.96 ;
     RECT  241.54 375.8 246.34 395.74 ;
     RECT  242.5 228.38 246.82 235.72 ;
     RECT  243.74 92.3 247.3 92.5 ;
     RECT  246.82 235.52 247.3 235.72 ;
     RECT  246.34 253.58 247.78 265.96 ;
     RECT  246.14 363.62 247.78 366.34 ;
     RECT  244.22 196.88 248.26 197.08 ;
     RECT  244.22 307.34 248.26 336.52 ;
     RECT  248.26 307.34 248.54 335.68 ;
     RECT  247.78 253.58 248.74 257.14 ;
     RECT  247.78 265.76 249.22 265.96 ;
     RECT  246.34 375.8 249.22 376 ;
     RECT  248.54 306.5 249.7 335.68 ;
     RECT  242.5 130.94 250.18 131.14 ;
     RECT  249.7 311.54 250.18 335.68 ;
     RECT  237.98 149.42 250.46 150.88 ;
     RECT  241.54 179.66 250.66 179.86 ;
     RECT  248.74 256.1 250.66 257.14 ;
     RECT  250.18 329.18 250.66 335.68 ;
     RECT  250.46 149.42 250.94 151.3 ;
     RECT  250.66 256.1 251.14 256.72 ;
     RECT  250.18 311.54 251.62 318.04 ;
     RECT  250.66 334.22 251.62 335.68 ;
     RECT  233.66 69.2 252.1 69.4 ;
     RECT  250.94 143.54 252.1 153.4 ;
     RECT  251.62 311.54 252.1 317.62 ;
     RECT  247.78 366.14 252.38 366.34 ;
     RECT  243.26 111.2 252.58 115.6 ;
     RECT  252.1 143.54 252.58 150.88 ;
     RECT  252.1 311.54 252.58 317.2 ;
     RECT  252.58 114.98 254.3 115.6 ;
     RECT  253.34 125.06 254.3 125.26 ;
     RECT  251.9 201.08 254.3 201.28 ;
     RECT  253.82 270.38 254.3 270.58 ;
     RECT  243.46 279.2 254.3 293.68 ;
     RECT  254.3 201.08 254.5 203.8 ;
     RECT  242.78 348.5 254.78 348.7 ;
     RECT  254.78 348.5 255.26 351.64 ;
     RECT  255.26 345.56 256.42 351.64 ;
     RECT  253.34 213.26 256.7 213.46 ;
     RECT  252.38 366.14 256.7 372.22 ;
     RECT  252.58 315.74 256.9 315.94 ;
     RECT  254.78 141.44 258.82 141.64 ;
     RECT  254.5 203.6 259.1 203.8 ;
     RECT  256.7 213.26 259.1 215.98 ;
     RECT  254.3 114.98 259.58 125.26 ;
     RECT  251.62 335.48 259.78 335.68 ;
     RECT  257.66 175.46 260.54 175.66 ;
     RECT  252.38 186.38 260.54 186.58 ;
     RECT  254.3 270.38 260.54 293.68 ;
     RECT  260.06 240.98 261.02 241.18 ;
     RECT  260.54 175.46 261.7 186.58 ;
     RECT  261.02 235.94 261.7 241.18 ;
     RECT  261.7 175.46 261.98 180.28 ;
     RECT  260.54 270.38 261.98 295.78 ;
     RECT  258.14 253.58 262.46 253.78 ;
     RECT  256.7 365.3 262.94 372.22 ;
     RECT  262.46 252.32 263.42 253.78 ;
     RECT  261.98 167.9 263.9 180.28 ;
     RECT  263.42 252.32 264.86 254.62 ;
     RECT  261.98 268.28 264.86 295.78 ;
     RECT  246.34 390.92 264.86 395.74 ;
     RECT  264.86 252.32 266.02 295.78 ;
     RECT  256.42 345.56 266.02 349.96 ;
     RECT  259.1 203.6 266.78 215.98 ;
     RECT  262.46 190.58 267.26 190.78 ;
     RECT  266.78 203.6 267.26 216.82 ;
     RECT  256.7 226.7 267.26 226.9 ;
     RECT  261.7 235.94 267.26 236.14 ;
     RECT  264.86 387.14 267.46 395.74 ;
     RECT  262.94 363.2 267.74 372.22 ;
     RECT  267.26 190.58 267.94 216.82 ;
     RECT  267.94 190.58 268.42 215.56 ;
     RECT  267.46 390.92 268.42 395.74 ;
     RECT  267.74 361.1 269.66 372.22 ;
     RECT  255.74 99.44 270.14 99.64 ;
     RECT  259.58 114.98 270.14 126.94 ;
     RECT  268.42 190.58 270.34 213.46 ;
     RECT  267.26 226.7 271.1 236.14 ;
     RECT  268.42 391.34 271.3 395.74 ;
     RECT  270.34 190.58 273.22 209.68 ;
     RECT  269.66 309.02 273.22 309.22 ;
     RECT  271.1 226.7 273.5 243.28 ;
     RECT  273.5 226.7 273.7 243.7 ;
     RECT  252.58 150.68 273.98 150.88 ;
     RECT  263.9 164.54 273.98 180.28 ;
     RECT  266.02 345.56 274.46 349.54 ;
     RECT  269.66 361.1 274.46 376.42 ;
     RECT  270.14 99.44 275.42 126.94 ;
     RECT  265.34 136.82 275.42 137.02 ;
     RECT  273.98 150.68 275.62 180.28 ;
     RECT  273.22 190.58 276.58 203.8 ;
     RECT  266.02 252.32 277.34 255.88 ;
     RECT  266.02 266.18 277.34 295.78 ;
     RECT  277.34 252.32 278.02 295.78 ;
     RECT  183.94 409.4 278.3 409.6 ;
     RECT  278.3 408.98 278.5 409.6 ;
     RECT  275.42 99.44 278.78 137.02 ;
     RECT  275.62 150.68 278.98 173.56 ;
     RECT  276.58 190.58 278.98 198.76 ;
     RECT  278.02 275.84 278.98 295.78 ;
     RECT  278.02 252.32 280.42 267.22 ;
     RECT  278.78 99.44 281.38 141.22 ;
     RECT  278.98 191 281.38 198.76 ;
     RECT  278.98 156.98 281.86 173.56 ;
     RECT  274.46 345.56 282.34 376.42 ;
     RECT  282.34 345.56 282.82 368.86 ;
     RECT  271.58 70.04 284.26 70.24 ;
     RECT  282.82 348.5 284.26 368.86 ;
     RECT  281.38 99.44 284.74 135.34 ;
     RECT  280.42 252.32 285.22 256.3 ;
     RECT  280.42 266.18 285.22 267.22 ;
     RECT  284.74 99.44 285.5 125.68 ;
     RECT  271.3 395.54 285.7 395.74 ;
     RECT  285.5 95.66 286.66 125.68 ;
     RECT  278.98 277.52 287.42 295.78 ;
     RECT  281.86 156.98 288.86 157.18 ;
     RECT  288.38 209.48 288.86 209.68 ;
     RECT  285.22 252.32 289.54 255.46 ;
     RECT  273.7 226.7 289.82 236.14 ;
     RECT  284.26 354.38 290.5 368.86 ;
     RECT  277.34 81.38 290.78 81.58 ;
     RECT  281.38 191 290.98 196.24 ;
     RECT  288.86 207.8 290.98 209.68 ;
     RECT  289.54 252.32 290.98 254.62 ;
     RECT  287.42 274.16 291.94 295.78 ;
     RECT  283.1 322.88 292.22 330.64 ;
     RECT  288.86 149.42 292.9 157.18 ;
     RECT  290.5 368.24 293.18 368.86 ;
     RECT  289.82 226.7 293.38 238.24 ;
     RECT  291.94 274.16 293.38 288.64 ;
     RECT  290.78 81.38 293.86 82 ;
     RECT  286.66 107.42 294.34 125.68 ;
     RECT  286.66 95.66 294.82 95.86 ;
     RECT  292.9 153.2 294.82 157.18 ;
     RECT  284.74 134.3 295.1 135.34 ;
     RECT  292.22 318.26 295.3 330.64 ;
     RECT  290.98 252.32 295.78 253.78 ;
     RECT  294.34 114.98 296.26 125.68 ;
     RECT  295.1 134.3 296.54 137.44 ;
     RECT  296.54 134.3 296.74 137.86 ;
     RECT  293.38 226.7 296.74 235.72 ;
     RECT  296.26 114.98 297.22 125.26 ;
     RECT  293.38 274.16 297.22 285.28 ;
     RECT  294.82 156.98 297.7 157.18 ;
     RECT  293.18 368.24 297.7 369.28 ;
     RECT  295.78 253.58 298.18 253.78 ;
     RECT  295.3 318.26 298.46 326.86 ;
     RECT  295.1 308.18 298.94 308.38 ;
     RECT  293.86 81.8 299.14 82 ;
     RECT  296.74 136.82 299.62 137.86 ;
     RECT  298.46 317.84 300.1 326.86 ;
     RECT  290.5 354.38 300.1 359.62 ;
     RECT  299.62 136.82 301.06 137.02 ;
     RECT  297.7 369.08 301.06 369.28 ;
     RECT  300.1 354.38 301.54 354.58 ;
     RECT  297.22 276.26 301.82 285.28 ;
     RECT  296.54 92.72 302.02 92.92 ;
     RECT  298.94 305.66 302.02 308.38 ;
     RECT  281.86 166.64 302.3 173.56 ;
     RECT  290.98 196.04 302.3 196.24 ;
     RECT  290.98 207.8 302.3 208 ;
     RECT  300.1 317.84 302.3 320.56 ;
     RECT  302.3 166.64 302.5 173.98 ;
     RECT  296.74 226.7 302.5 226.9 ;
     RECT  301.82 276.26 302.5 287.38 ;
     RECT  297.5 337.58 302.5 337.78 ;
     RECT  302.3 196.04 302.78 208 ;
     RECT  302.3 239.72 302.78 239.92 ;
     RECT  302.5 276.26 303.46 278.14 ;
     RECT  302.5 287.18 303.46 287.38 ;
     RECT  302.3 380 303.46 380.2 ;
     RECT  302.78 239.72 304.42 241.18 ;
     RECT  303.26 217.04 304.9 217.24 ;
     RECT  302.5 173.78 305.66 173.98 ;
     RECT  301.34 182.6 305.66 182.8 ;
     RECT  304.42 239.72 305.66 239.92 ;
     RECT  302.3 257.78 306.14 257.98 ;
     RECT  297.22 114.98 307.1 122.74 ;
     RECT  306.14 257.78 307.3 263.44 ;
     RECT  303.74 290.54 307.78 290.74 ;
     RECT  302.3 311.96 308.54 320.56 ;
     RECT  307.58 330.02 308.54 330.22 ;
     RECT  302.78 194.78 309.5 208 ;
     RECT  305.66 233 310.94 239.92 ;
     RECT  309.02 360.26 311.42 360.46 ;
     RECT  303.46 277.1 311.9 278.14 ;
     RECT  309.5 194.78 312.58 208.84 ;
     RECT  311.9 273.74 312.86 278.14 ;
     RECT  308.06 219.56 314.02 219.76 ;
     RECT  308.06 248.96 314.02 249.16 ;
     RECT  311.42 355.22 314.3 360.46 ;
     RECT  312.58 194.78 314.5 205.9 ;
     RECT  307.3 257.78 315.26 257.98 ;
     RECT  314.3 355.22 316.7 361.3 ;
     RECT  308.54 311.96 317.18 330.22 ;
     RECT  317.18 311.12 317.38 330.22 ;
     RECT  305.66 173.78 317.66 182.8 ;
     RECT  314.5 194.78 317.66 205.48 ;
     RECT  315.26 251.9 317.66 257.98 ;
     RECT  316.7 355.22 318.34 362.56 ;
     RECT  307.1 114.98 318.62 130.3 ;
     RECT  312.86 273.74 318.62 285.28 ;
     RECT  317.38 311.12 318.62 323.5 ;
     RECT  310.94 228.38 319.58 239.92 ;
     RECT  318.34 355.22 320.06 361.3 ;
     RECT  318.62 272.9 320.26 286.12 ;
     RECT  319.58 223.76 320.74 239.92 ;
     RECT  320.06 349.76 321.22 361.3 ;
     RECT  320.26 273.74 321.5 286.12 ;
     RECT  320.74 230.9 321.7 239.92 ;
     RECT  321.7 231.32 322.18 239.92 ;
     RECT  317.66 251.9 322.66 260.92 ;
     RECT  317.66 173.78 323.62 205.48 ;
     RECT  321.22 361.1 323.62 361.3 ;
     RECT  318.62 114.98 323.9 134.5 ;
     RECT  323.9 111.62 324.1 134.5 ;
     RECT  323.62 173.78 326.02 173.98 ;
     RECT  323.62 182.6 326.02 205.48 ;
     RECT  322.18 232.58 326.78 239.92 ;
     RECT  322.66 251.9 326.78 256.72 ;
     RECT  324.1 111.62 327.26 130.3 ;
     RECT  318.62 303.98 327.46 323.5 ;
     RECT  329.18 145.22 330.62 145.42 ;
     RECT  323.42 164.12 330.82 164.32 ;
     RECT  321.22 349.76 331.1 349.96 ;
     RECT  321.5 273.74 331.3 292.84 ;
     RECT  325.82 338.42 331.58 338.62 ;
     RECT  326.78 232.58 332.06 256.72 ;
     RECT  331.3 273.74 333.22 278.14 ;
     RECT  331.58 331.28 333.22 338.62 ;
     RECT  331.1 349.76 333.22 350.38 ;
     RECT  330.62 145.22 333.98 153.4 ;
     RECT  327.26 107.42 334.66 130.3 ;
     RECT  326.02 182.6 334.94 202.54 ;
     RECT  334.66 118.76 336.1 130.3 ;
     RECT  327.46 303.98 336.1 317.2 ;
     RECT  336.1 119.6 336.58 130.3 ;
     RECT  331.3 292.64 336.58 292.84 ;
     RECT  334.94 368.24 337.54 368.44 ;
     RECT  333.98 141.44 338.02 153.4 ;
     RECT  332.06 232.58 338.3 260.08 ;
     RECT  334.94 182.6 338.5 215.98 ;
     RECT  333.22 338.42 338.5 338.62 ;
     RECT  338.5 182.6 339.94 210.1 ;
     RECT  339.94 194.78 340.42 210.1 ;
     RECT  333.22 277.52 341.18 278.14 ;
     RECT  340.42 194.78 341.38 209.68 ;
     RECT  341.18 277.52 341.38 281.92 ;
     RECT  338.3 229.22 341.66 260.08 ;
     RECT  341.66 228.8 343.58 260.08 ;
     RECT  339.94 182.6 343.78 183.22 ;
     RECT  343.58 228.38 343.78 260.08 ;
     RECT  333.22 349.76 345.02 349.96 ;
     RECT  336.58 126.32 346.94 130.3 ;
     RECT  338.02 141.44 346.94 145.42 ;
     RECT  341.38 194.78 347.14 205.9 ;
     RECT  346.94 126.32 347.62 145.42 ;
     RECT  336.86 103.64 348.1 103.84 ;
     RECT  343.78 228.38 348.1 243.28 ;
     RECT  345.02 345.98 348.1 349.96 ;
     RECT  347.14 202.34 348.58 205.9 ;
     RECT  343.78 256.1 348.58 260.08 ;
     RECT  348.1 228.8 349.06 237.82 ;
     RECT  348.1 345.98 349.06 346.18 ;
     RECT  343.78 183.02 350.5 183.22 ;
     RECT  348.58 205.7 350.5 205.9 ;
     RECT  342.14 70.04 351.94 70.24 ;
     RECT  349.06 229.22 351.94 237.82 ;
     RECT  341.38 277.52 352.7 281.5 ;
     RECT  336.1 308.18 352.7 317.2 ;
     RECT  347.62 133.46 352.9 137.44 ;
     RECT  348.58 256.1 352.9 256.3 ;
     RECT  352.7 164.12 353.66 164.32 ;
     RECT  352.7 277.52 353.66 289.06 ;
     RECT  353.66 275 354.62 289.06 ;
     RECT  352.9 133.46 356.06 133.66 ;
     RECT  354.62 272.9 357.02 289.06 ;
     RECT  357.02 272.48 357.98 289.06 ;
     RECT  356.06 125.06 358.46 133.66 ;
     RECT  352.7 305.66 359.42 317.2 ;
     RECT  353.66 164.12 359.62 171.46 ;
     RECT  359.42 345.98 360.86 346.18 ;
     RECT  357.98 266.6 361.34 289.06 ;
     RECT  359.42 305.66 361.34 319.3 ;
     RECT  361.34 304.4 363.74 319.3 ;
     RECT  358.46 122.54 363.94 133.66 ;
     RECT  361.34 266.18 364.22 289.06 ;
     RECT  363.74 303.14 364.22 319.3 ;
     RECT  359.62 166.22 364.7 171.46 ;
     RECT  363.94 122.54 366.34 130.72 ;
     RECT  351.94 237.62 368.06 237.82 ;
     RECT  364.7 166.22 368.74 172.3 ;
     RECT  366.14 100.28 369.22 100.48 ;
     RECT  368.06 235.1 369.7 237.82 ;
     RECT  369.7 235.52 369.98 237.82 ;
     RECT  368.74 172.1 371.14 172.3 ;
     RECT  369.98 254.84 371.14 255.04 ;
     RECT  364.22 266.18 371.14 319.3 ;
     RECT  368.06 334.22 371.62 334.42 ;
     RECT  361.82 145.64 372.58 145.84 ;
     RECT  369.98 235.52 372.58 244.12 ;
     RECT  371.14 272.48 372.86 319.3 ;
     RECT  359.42 186.8 373.34 187 ;
     RECT  372.86 272.48 374.3 319.72 ;
     RECT  365.18 201.08 374.5 201.28 ;
     RECT  366.34 129.68 375.74 130.72 ;
     RECT  374.3 272.48 377.18 322.66 ;
     RECT  360.86 345.98 377.18 350.38 ;
     RECT  377.18 272.48 377.38 327.28 ;
     RECT  378.14 262.82 379.58 263.02 ;
     RECT  375.74 129.26 379.78 130.72 ;
     RECT  377.38 272.48 379.78 289.06 ;
     RECT  377.38 303.98 379.78 327.28 ;
     RECT  377.18 341.78 379.78 350.38 ;
     RECT  379.58 255.26 380.06 263.02 ;
     RECT  379.78 272.48 380.06 286.54 ;
     RECT  373.34 180.5 380.26 187 ;
     RECT  372.58 235.52 381.02 241.18 ;
     RECT  380.06 255.26 381.02 286.54 ;
     RECT  381.02 235.1 381.22 241.18 ;
     RECT  369.5 77.6 382.18 77.8 ;
     RECT  371.42 104.06 382.18 111.82 ;
     RECT  381.22 235.52 382.18 241.18 ;
     RECT  380.26 180.5 382.66 180.7 ;
     RECT  380.54 191 382.66 191.2 ;
     RECT  381.02 251.06 383.14 286.54 ;
     RECT  379.78 303.98 383.14 323.5 ;
     RECT  379.78 341.78 383.14 349.96 ;
     RECT  383.14 251.06 384.1 283.6 ;
     RECT  384.1 251.06 384.58 266.8 ;
     RECT  383.14 348.92 385.06 349.96 ;
     RECT  382.18 235.94 385.54 241.18 ;
     RECT  382.18 111.2 385.82 111.82 ;
     RECT  381.02 122.54 385.82 122.74 ;
     RECT  383.14 303.98 385.82 310.9 ;
     RECT  384.58 251.06 386.02 255.46 ;
     RECT  384.1 277.94 386.5 282.34 ;
     RECT  385.82 111.2 387.94 122.74 ;
     RECT  385.54 237.62 387.94 241.18 ;
     RECT  385.82 296.42 387.94 310.9 ;
     RECT  386.02 251.06 388.42 251.26 ;
     RECT  382.46 100.28 388.9 100.48 ;
     RECT  387.94 240.98 388.9 241.18 ;
     RECT  386.78 194.78 389.86 197.5 ;
     RECT  386.5 280.04 390.34 282.34 ;
     RECT  390.34 282.14 390.82 282.34 ;
     RECT  387.94 302.72 390.82 310.9 ;
     RECT  389.86 194.78 391.3 194.98 ;
     RECT  375.74 142.28 392.26 143.32 ;
     RECT  392.26 142.28 392.74 142.48 ;
     RECT  383.14 322.88 392.74 323.5 ;
     RECT  387.94 111.2 393.7 111.4 ;
     RECT  390.82 308.18 394.18 310.9 ;
     RECT  367.1 213.26 394.66 213.46 ;
     RECT  394.18 308.18 394.66 308.38 ;
     RECT  384.58 266.6 398.02 266.8 ;
     RECT  392.74 322.88 398.02 323.08 ;
     RECT  385.06 349.76 398.02 349.96 ;
     RECT  387.94 122.54 399.94 122.74 ;
     RECT  384.38 172.1 399.94 172.3 ;
  END
END cve2_register_file_ff
END LIBRARY
