module timer_unit (gnt_o,
    r_opc_o,
    busy_o,
    clk_i,
    event_hi_i,
    event_lo_i,
    irq_hi_o,
    irq_lo_o,
    r_valid_o,
    ref_clk_i,
    req_i,
    rst_ni,
    wen_i,
    addr_i,
    be_i,
    id_i,
    r_id_o,
    r_rdata_o,
    wdata_i);
 output gnt_o;
 output r_opc_o;
 output busy_o;
 input clk_i;
 input event_hi_i;
 input event_lo_i;
 output irq_hi_o;
 output irq_lo_o;
 output r_valid_o;
 input ref_clk_i;
 input req_i;
 input rst_ni;
 input wen_i;
 input [31:0] addr_i;
 input [3:0] be_i;
 input [4:0] id_i;
 output [4:0] r_id_o;
 output [31:0] r_rdata_o;
 input [31:0] wdata_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire net56;
 wire net55;
 wire _0233_;
 wire _0234_;
 wire net54;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire net53;
 wire net52;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire net51;
 wire net50;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire net49;
 wire _0262_;
 wire _0263_;
 wire net48;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire net47;
 wire net46;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire net45;
 wire net44;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire net43;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire net42;
 wire _0470_;
 wire net41;
 wire net40;
 wire _0473_;
 wire net39;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire net38;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire net37;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire net36;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire net35;
 wire net34;
 wire _0586_;
 wire net33;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire net32;
 wire net31;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire net30;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire net29;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire net28;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire net27;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire net26;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire net25;
 wire _0731_;
 wire net24;
 wire _0733_;
 wire _0734_;
 wire net23;
 wire _0736_;
 wire _0737_;
 wire net22;
 wire _0739_;
 wire net21;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire net20;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire net19;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire net18;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire net17;
 wire net16;
 wire _0796_;
 wire _0797_;
 wire net15;
 wire net14;
 wire _0800_;
 wire net13;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire net12;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire net11;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire net10;
 wire _0852_;
 wire _0853_;
 wire net9;
 wire net8;
 wire _0856_;
 wire net7;
 wire _0858_;
 wire _0859_;
 wire net6;
 wire _0861_;
 wire net5;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire net4;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire net3;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire net79;
 wire net78;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire net77;
 wire net76;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire net75;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire net74;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire net73;
 wire net72;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire net66;
 wire net65;
 wire _1031_;
 wire _1032_;
 wire net64;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire net63;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire net62;
 wire net61;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire net60;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire net59;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire net58;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire net57;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire net90;
 wire net2;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_10_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_10_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_11_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_11_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_12_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_12_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_13_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_13_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_14_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_14_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_1_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_1_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_2_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_2_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_3_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_3_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_4_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_4_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_5_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_5_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_6_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_6_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_7_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_7_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_8_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_8_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_9_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_9_B ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ;
 wire \counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ;
 wire \counter_hi_i.target_reached_o ;
 wire \counter_hi_i.target_reached_o_reg_D ;
 wire \counter_lo_i.enable_count_i_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_B ;
 wire \counter_lo_i.target_reached_o ;
 wire \counter_lo_i.target_reached_o_reg_D ;
 wire \prescaler_hi_i.enable_count_i_$_AND__Y_B_$_MUX__Y_S_$_AND__Y_B ;
 wire \prescaler_hi_i.target_reached_o ;
 wire \prescaler_hi_i.target_reached_o_$_MUX__A_S_$_AND__Y_A ;
 wire \prescaler_hi_i.target_reached_o_reg_D ;
 wire \prescaler_lo_i.target_reached_o ;
 wire \prescaler_lo_i.target_reached_o_reg_D ;
 wire \s_addr_$_NOT__A_1_Y ;
 wire \s_addr_$_NOT__A_2_Y ;
 wire \s_addr_$_NOT__A_Y ;
 wire \s_cfg_hi_$_OR__Y_A_$_MUX__Y_S_$_AND__Y_A_$_AND__Y_A ;
 wire s_ref_clk0;
 wire s_ref_clk1;
 wire s_ref_clk2;
 wire s_ref_clk3;
 wire \s_ref_clk_edge_$_AND__Y_B ;
 wire \s_ref_clk_edge_del_$_AND__Y_B ;
 wire \s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ;
 wire s_wen;
 wire VDD;
 wire VSS;
 wire net1;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_0_clk_i;
 wire clknet_3_0__leaf_clk_i;
 wire clknet_3_1__leaf_clk_i;
 wire clknet_3_2__leaf_clk_i;
 wire clknet_3_3__leaf_clk_i;
 wire clknet_3_4__leaf_clk_i;
 wire clknet_3_5__leaf_clk_i;
 wire clknet_3_6__leaf_clk_i;
 wire clknet_3_7__leaf_clk_i;
 wire net113;
 wire net114;
 wire net115;
 wire [31:0] \counter_hi_i.compare_value_i ;
 wire [31:0] \counter_hi_i.enable_count_i_$_MUX__S_31_B ;
 wire [0:0] \counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B ;
 wire [31:0] \counter_hi_i.s_count ;
 wire [31:0] \counter_lo_i.compare_value_i ;
 wire [31:0] \counter_lo_i.enable_count_i_$_MUX__S_31_B ;
 wire [0:0] \counter_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B ;
 wire [31:0] \counter_lo_i.s_count ;
 wire [7:0] \prescaler_hi_i.compare_value_i ;
 wire [31:0] \prescaler_hi_i.enable_count_i_$_MUX__S_31_B ;
 wire [0:0] \prescaler_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B ;
 wire [31:0] \prescaler_hi_i.s_count ;
 wire [7:0] \prescaler_lo_i.compare_value_i ;
 wire [31:0] \prescaler_lo_i.enable_count_i_$_MUX__S_31_B ;
 wire [0:0] \prescaler_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B ;
 wire [31:0] \prescaler_lo_i.s_count ;
 wire [5:0] s_addr;
 wire [5:0] s_cfg_hi;
 wire [31:0] s_cfg_hi_reg;
 wire [5:0] s_cfg_lo;
 wire [31:0] s_cfg_lo_reg;

 sg13g2_inv_1 _1449_ (.VDD(VDD),
    .Y(_0934_),
    .A(s_cfg_hi_reg[0]),
    .VSS(VSS));
 sg13g2_inv_1 _1450_ (.VDD(VDD),
    .Y(_0935_),
    .A(s_cfg_lo_reg[0]),
    .VSS(VSS));
 sg13g2_nand2_2 _1451_ (.Y(busy_o),
    .A(_0934_),
    .B(_0935_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1452_ (.VDD(VDD),
    .Y(_0936_),
    .A(addr_i[4]),
    .VSS(VSS));
 sg13g2_nand2b_1 _1453_ (.Y(_0937_),
    .B(req_i),
    .A_N(wen_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _1454_ (.A(_0936_),
    .B(addr_i[5]),
    .C(_0937_),
    .Y(_0938_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1455_ (.A(addr_i[0]),
    .B(addr_i[1]),
    .Y(_0939_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _1456_ (.A(addr_i[3]),
    .B_N(addr_i[2]),
    .Y(_0940_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _1457_ (.A(_0939_),
    .B(_0940_),
    .X(_0941_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _1458_ (.A(_0938_),
    .B(_0941_),
    .X(_0942_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net92),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(net92),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1461_ (.A0(\counter_hi_i.compare_value_i [0]),
    .A1(wdata_i[0]),
    .S(net109),
    .X(_0000_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1462_ (.A0(\counter_hi_i.compare_value_i [10]),
    .A1(wdata_i[10]),
    .S(net111),
    .X(_0001_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1463_ (.A0(\counter_hi_i.compare_value_i [11]),
    .A1(wdata_i[11]),
    .S(net110),
    .X(_0002_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1464_ (.A0(\counter_hi_i.compare_value_i [12]),
    .A1(wdata_i[12]),
    .S(net110),
    .X(_0003_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1465_ (.A0(\counter_hi_i.compare_value_i [13]),
    .A1(wdata_i[13]),
    .S(net110),
    .X(_0004_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1466_ (.A0(\counter_hi_i.compare_value_i [14]),
    .A1(wdata_i[14]),
    .S(net110),
    .X(_0005_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1467_ (.A0(\counter_hi_i.compare_value_i [15]),
    .A1(wdata_i[15]),
    .S(net108),
    .X(_0006_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1468_ (.A0(\counter_hi_i.compare_value_i [16]),
    .A1(wdata_i[16]),
    .S(net109),
    .X(_0007_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout87 (.A(_0468_),
    .X(net87),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1470_ (.A0(\counter_hi_i.compare_value_i [17]),
    .A1(wdata_i[17]),
    .S(net108),
    .X(_0008_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1471_ (.A0(\counter_hi_i.compare_value_i [18]),
    .A1(wdata_i[18]),
    .S(net108),
    .X(_0009_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(net87),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1473_ (.A0(\counter_hi_i.compare_value_i [19]),
    .A1(wdata_i[19]),
    .S(net108),
    .X(_0010_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1474_ (.A0(\counter_hi_i.compare_value_i [1]),
    .A1(wdata_i[1]),
    .S(net109),
    .X(_0011_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1475_ (.A0(\counter_hi_i.compare_value_i [20]),
    .A1(wdata_i[20]),
    .S(net108),
    .X(_0012_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1476_ (.A0(\counter_hi_i.compare_value_i [21]),
    .A1(wdata_i[21]),
    .S(net107),
    .X(_0013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout85 (.A(net87),
    .X(net85),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1478_ (.A0(\counter_hi_i.compare_value_i [22]),
    .A1(wdata_i[22]),
    .S(net107),
    .X(_0014_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1479_ (.A0(\counter_hi_i.compare_value_i [23]),
    .A1(wdata_i[23]),
    .S(net107),
    .X(_0015_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net87),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1481_ (.A0(\counter_hi_i.compare_value_i [24]),
    .A1(wdata_i[24]),
    .S(net108),
    .X(_0016_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1482_ (.A0(\counter_hi_i.compare_value_i [25]),
    .A1(wdata_i[25]),
    .S(net107),
    .X(_0017_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_0468_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1484_ (.A0(\counter_hi_i.compare_value_i [26]),
    .A1(wdata_i[26]),
    .S(net108),
    .X(_0018_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1485_ (.A0(\counter_hi_i.compare_value_i [27]),
    .A1(wdata_i[27]),
    .S(net107),
    .X(_0019_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_0468_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1487_ (.A0(\counter_hi_i.compare_value_i [28]),
    .A1(wdata_i[28]),
    .S(net107),
    .X(_0020_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1488_ (.A0(\counter_hi_i.compare_value_i [29]),
    .A1(wdata_i[29]),
    .S(net107),
    .X(_0021_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1489_ (.A0(\counter_hi_i.compare_value_i [2]),
    .A1(wdata_i[2]),
    .S(net109),
    .X(_0022_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1490_ (.A0(\counter_hi_i.compare_value_i [30]),
    .A1(wdata_i[30]),
    .S(net107),
    .X(_0023_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1491_ (.A0(\counter_hi_i.compare_value_i [31]),
    .A1(wdata_i[31]),
    .S(net109),
    .X(_0024_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1492_ (.A0(\counter_hi_i.compare_value_i [3]),
    .A1(wdata_i[3]),
    .S(net110),
    .X(_0025_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1493_ (.A0(\counter_hi_i.compare_value_i [4]),
    .A1(wdata_i[4]),
    .S(net109),
    .X(_0026_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1494_ (.A0(\counter_hi_i.compare_value_i [5]),
    .A1(wdata_i[5]),
    .S(net109),
    .X(_0027_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1495_ (.A0(\counter_hi_i.compare_value_i [6]),
    .A1(wdata_i[6]),
    .S(net109),
    .X(_0028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1496_ (.A0(\counter_hi_i.compare_value_i [7]),
    .A1(wdata_i[7]),
    .S(net111),
    .X(_0029_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1497_ (.A0(\counter_hi_i.compare_value_i [8]),
    .A1(wdata_i[8]),
    .S(net110),
    .X(_0030_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout81 (.A(_0473_),
    .X(net81),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1500_ (.A0(\counter_hi_i.compare_value_i [9]),
    .A1(wdata_i[9]),
    .S(net110),
    .X(_0031_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1501_ (.VDD(VDD),
    .Y(_0953_),
    .A(s_cfg_hi_reg[1]),
    .VSS(VSS));
 sg13g2_nor2b_1 _1502_ (.A(s_cfg_lo_reg[31]),
    .B_N(s_cfg_hi_reg[4]),
    .Y(_0954_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _1503_ (.X(_0955_),
    .A(s_cfg_lo_reg[31]),
    .B(s_cfg_lo_reg[4]),
    .C(\counter_lo_i.target_reached_o ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1504_ (.B1(\counter_hi_i.target_reached_o ),
    .VDD(VDD),
    .Y(_0956_),
    .VSS(VSS),
    .A1(_0954_),
    .A2(_0955_));
 sg13g2_nor2b_1 _1505_ (.A(wen_i),
    .B_N(req_i),
    .Y(_0957_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _1506_ (.A(addr_i[4]),
    .B_N(addr_i[5]),
    .Y(_0958_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1507_ (.B(_0939_),
    .C(_0940_),
    .A(_0957_),
    .Y(_0959_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0958_));
 sg13g2_and3_1 _1508_ (.X(_0960_),
    .A(_0953_),
    .B(_0956_),
    .C(_0959_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout79 (.A(net81),
    .X(net79),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout78 (.A(_0473_),
    .X(net78),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1511_ (.VDD(VDD),
    .Y(_0963_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .VSS(VSS));
 sg13g2_nand3_1 _1512_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .Y(_0964_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1513_ (.VDD(VDD),
    .Y(_0965_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .VSS(VSS));
 sg13g2_buf_2 fanout77 (.A(net78),
    .X(net77),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(_1028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1516_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .Y(_0968_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _1517_ (.A(_0965_),
    .B(_0968_),
    .Y(_0969_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1518_ (.Y(_0970_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .B(_0969_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 _1520_ (.X(_0972_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1521_ (.B(net112),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .Y(_0973_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0972_));
 sg13g2_nand2_1 _1522_ (.Y(_0974_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 _1523_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0975_),
    .B(_0974_),
    .A(_0973_));
 sg13g2_or4_2 _1524_ (.A(_0963_),
    .B(_0964_),
    .C(_0970_),
    .D(_0975_),
    .X(_0976_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _1525_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0977_),
    .B(\prescaler_hi_i.target_reached_o ),
    .A(s_cfg_hi_reg[7]));
 sg13g2_nand2_2 _1526_ (.Y(_0978_),
    .A(s_ref_clk1),
    .B(\s_ref_clk_edge_$_AND__Y_B ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1527_ (.B(\prescaler_hi_i.target_reached_o_$_MUX__A_S_$_AND__Y_A ),
    .C(_0978_),
    .A(s_cfg_hi_reg[7]),
    .Y(_0979_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _1528_ (.A2(_0979_),
    .A1(_0977_),
    .B1(\prescaler_hi_i.enable_count_i_$_AND__Y_B_$_MUX__Y_S_$_AND__Y_B ),
    .X(_0980_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1529_ (.B1(s_cfg_hi_reg[0]),
    .VDD(VDD),
    .Y(_0981_),
    .VSS(VSS),
    .A1(\prescaler_hi_i.target_reached_o_$_MUX__A_S_$_AND__Y_A ),
    .A2(\prescaler_hi_i.target_reached_o ));
 sg13g2_a21oi_1 _1530_ (.VSS(VSS),
    .VDD(VDD),
    .A1(s_cfg_lo_reg[0]),
    .A2(s_cfg_lo_reg[31]),
    .Y(_0982_),
    .B1(_0981_));
 sg13g2_nand2b_1 _1531_ (.Y(_0983_),
    .B(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ),
    .A_N(\counter_lo_i.enable_count_i_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_B ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _1532_ (.Y(_0984_),
    .B(s_cfg_lo_reg[6]),
    .A_N(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1533_ (.VDD(VDD),
    .Y(_0985_),
    .A(s_cfg_lo_reg[7]),
    .VSS(VSS));
 sg13g2_a221oi_1 _1534_ (.VSS(VSS),
    .VDD(VDD),
    .B2(_0984_),
    .C1(_0985_),
    .B1(_0983_),
    .A1(s_ref_clk2),
    .Y(_0986_),
    .A2(\s_ref_clk_edge_del_$_AND__Y_B ));
 sg13g2_nor2_1 _1535_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_12_B ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_2_A ),
    .Y(_0987_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1536_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_14_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_14_B ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_A ),
    .D(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_B ),
    .Y(_0988_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1537_ (.Y(_0989_),
    .A(_0987_),
    .B(_0988_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1538_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_10_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_10_B ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_11_A ),
    .D(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_11_B ),
    .Y(_0990_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1539_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_12_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_13_A ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_13_B ),
    .D(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_2_B ),
    .Y(_0991_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1540_ (.Y(_0992_),
    .A(_0990_),
    .B(_0991_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1541_ (.VDD(VDD),
    .Y(_0993_),
    .A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_7_A ),
    .VSS(VSS));
 sg13g2_nor2_1 _1542_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_9_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_9_B ),
    .Y(_0994_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _1543_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_1_A ),
    .Y(_0995_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_1_B ));
 sg13g2_nand4_1 _1544_ (.B(s_cfg_lo_reg[31]),
    .C(_0994_),
    .A(_0993_),
    .Y(_0996_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0995_));
 sg13g2_nor4_1 _1545_ (.A(_0986_),
    .B(_0989_),
    .C(_0992_),
    .D(_0996_),
    .Y(_0997_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1546_ (.VDD(VDD),
    .Y(_0998_),
    .A(\prescaler_lo_i.target_reached_o ),
    .VSS(VSS));
 sg13g2_o21ai_1 _1547_ (.B1(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ),
    .VDD(VDD),
    .Y(_0999_),
    .VSS(VSS),
    .A1(\counter_lo_i.enable_count_i_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_B ),
    .A2(s_cfg_lo_reg[7]));
 sg13g2_a21oi_2 _1548_ (.VSS(VSS),
    .VDD(VDD),
    .B1(_0935_),
    .Y(_1000_),
    .A2(_0999_),
    .A1(_0998_));
 sg13g2_nor3_1 _1549_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_3_B ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_4_A ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_4_B ),
    .Y(_1001_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1550_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_5_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_5_B ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_6_A ),
    .D(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_6_B ),
    .Y(_1002_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1551_ (.A(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_3_A ),
    .B(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_7_B ),
    .C(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_8_A ),
    .D(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_8_B ),
    .Y(_1003_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _1552_ (.A(_1000_),
    .B(_1001_),
    .C(_1002_),
    .D(_1003_),
    .X(_1004_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _1553_ (.Y(_1005_),
    .B1(_0997_),
    .B2(_1004_),
    .A2(_0982_),
    .A1(_0980_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(net76),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1555_ (.VDD(VDD),
    .Y(_1007_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .VSS(VSS));
 sg13g2_nand4_1 _1556_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .Y(_1008_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]));
 sg13g2_or2_1 _1557_ (.VSS(VSS),
    .VDD(VDD),
    .X(_1009_),
    .B(_1008_),
    .A(_1007_));
 sg13g2_buf_2 fanout73 (.A(_0242_),
    .X(net73),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _1560_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .X(_1012_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _1561_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .D(_1012_),
    .X(_1013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1562_ (.Y(_1014_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .B(_1013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _1563_ (.A(_0976_),
    .B(net28),
    .C(net106),
    .Y(_1015_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_1014_));
 sg13g2_nand4_1 _1564_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .Y(_1016_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_1015_));
 sg13g2_xor2_1 _1565_ (.B(_1016_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .X(_1017_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_2 _1566_ (.A(addr_i[4]),
    .B(addr_i[5]),
    .C(_0937_),
    .X(_1018_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1567_ (.B(addr_i[3]),
    .C(_0939_),
    .A(addr_i[2]),
    .Y(_1019_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _1568_ (.VSS(VSS),
    .VDD(VDD),
    .X(_1020_),
    .B(_1019_),
    .A(_1018_));
 sg13g2_buf_2 fanout71 (.A(_0242_),
    .X(net71),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout70 (.A(net71),
    .X(net70),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout69 (.A(net71),
    .X(net69),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout68 (.A(_0247_),
    .X(net68),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout67 (.A(_0247_),
    .X(net67),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1574_ (.A(wdata_i[31]),
    .B(net14),
    .Y(_1026_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1575_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1017_),
    .A2(net16),
    .Y(_1027_),
    .B1(_1026_));
 sg13g2_and2_1 _1576_ (.A(net7),
    .B(_1027_),
    .X(\counter_hi_i.s_count [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1577_ (.B(_0956_),
    .C(_0959_),
    .A(_0953_),
    .Y(_1028_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout66 (.A(_0247_),
    .X(net66),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1580_ (.A(wdata_i[30]),
    .B(net15),
    .Y(_1031_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1581_ (.A(_1018_),
    .B(_1019_),
    .Y(_1032_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout64 (.A(net66),
    .X(net64),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1583_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .C(_1015_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .Y(_1034_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1584_ (.Y(_1035_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .B(_1034_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1585_ (.A(net103),
    .B(_1035_),
    .Y(_1036_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1586_ (.A(net74),
    .B(_1031_),
    .C(_1036_),
    .Y(\counter_hi_i.s_count [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout63 (.A(_0589_),
    .X(net63),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _1588_ (.A(_0970_),
    .B(_0975_),
    .C(net28),
    .Y(_1038_),
    .VDD(VDD),
    .VSS(VSS),
    .D(net106));
 sg13g2_nand2b_1 _1589_ (.Y(_1039_),
    .B(_1038_),
    .A_N(_0964_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1590_ (.Y(_1040_),
    .A(_0963_),
    .B(_1039_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1591_ (.A(wdata_i[21]),
    .B(_1018_),
    .C(_1019_),
    .Y(_1041_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _1592_ (.Y(_1042_),
    .B(net8),
    .A_N(_1041_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1593_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net17),
    .A2(_1040_),
    .Y(\counter_hi_i.s_count [21]),
    .B1(_1042_));
 sg13g2_nor2_1 _1594_ (.A(wdata_i[20]),
    .B(net14),
    .Y(_1043_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1595_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .C(_1038_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .Y(_1044_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1596_ (.Y(_1045_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(_1044_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1597_ (.A(net104),
    .B(_1045_),
    .Y(_1046_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1598_ (.A(net76),
    .B(_1043_),
    .C(_1046_),
    .Y(\counter_hi_i.s_count [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _1599_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .B(_1038_),
    .X(_1047_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1600_ (.Y(_1048_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .B(_1047_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout62 (.A(net63),
    .X(net62),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout61 (.A(net63),
    .X(net61),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1603_ (.B1(net9),
    .VDD(VDD),
    .Y(_1051_),
    .VSS(VSS),
    .A1(wdata_i[19]),
    .A2(net12));
 sg13g2_a21oi_1 _1604_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net17),
    .A2(_1048_),
    .Y(\counter_hi_i.s_count [19]),
    .B1(_1051_));
 sg13g2_xnor2_1 _1605_ (.Y(_1052_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .B(_1038_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1606_ (.B1(net9),
    .VDD(VDD),
    .Y(_1053_),
    .VSS(VSS),
    .A1(wdata_i[18]),
    .A2(net11));
 sg13g2_a21oi_1 _1607_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net17),
    .A2(_1052_),
    .Y(\counter_hi_i.s_count [18]),
    .B1(_1053_));
 sg13g2_buf_2 fanout60 (.A(net63),
    .X(net60),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _1609_ (.A(_0975_),
    .B(net28),
    .C(net106),
    .Y(_1055_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _1610_ (.A(_0969_),
    .B(_1055_),
    .X(_1056_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1611_ (.Y(_1057_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .B(_1056_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1612_ (.B1(net8),
    .VDD(VDD),
    .Y(_1058_),
    .VSS(VSS),
    .A1(wdata_i[17]),
    .A2(net11));
 sg13g2_a21oi_1 _1613_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1057_),
    .Y(\counter_hi_i.s_count [17]),
    .B1(_1058_));
 sg13g2_nor2_1 _1614_ (.A(wdata_i[16]),
    .B(net14),
    .Y(_1059_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1615_ (.A(_0968_),
    .B(_0975_),
    .C(net28),
    .D(net106),
    .Y(_1060_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1616_ (.Y(_1061_),
    .A(_0965_),
    .B(_1060_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1617_ (.A(_1032_),
    .B(_1061_),
    .Y(_1062_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1618_ (.A(net76),
    .B(_1059_),
    .C(_1062_),
    .Y(\counter_hi_i.s_count [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1619_ (.Y(_1063_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1620_ (.A(_0973_),
    .B(_0974_),
    .Y(_1064_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _1621_ (.A(net28),
    .B(net106),
    .Y(_1065_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1622_ (.Y(_1066_),
    .A(_1064_),
    .B(_1065_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1623_ (.A(_1063_),
    .B(_1066_),
    .Y(_1067_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1624_ (.Y(_1068_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .B(_1067_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1625_ (.B1(net8),
    .VDD(VDD),
    .Y(_1069_),
    .VSS(VSS),
    .A1(wdata_i[15]),
    .A2(net11));
 sg13g2_a21oi_1 _1626_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1068_),
    .Y(\counter_hi_i.s_count [15]),
    .B1(_1069_));
 sg13g2_and3_1 _1627_ (.X(_1070_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .B(_1064_),
    .C(_1065_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1628_ (.Y(_1071_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .B(_1070_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1629_ (.B1(net9),
    .VDD(VDD),
    .Y(_1072_),
    .VSS(VSS),
    .A1(wdata_i[14]),
    .A2(net12));
 sg13g2_a21oi_1 _1630_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1071_),
    .Y(\counter_hi_i.s_count [14]),
    .B1(_1072_));
 sg13g2_xnor2_1 _1631_ (.Y(_1073_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .B(_1055_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1632_ (.B1(net8),
    .VDD(VDD),
    .Y(_1074_),
    .VSS(VSS),
    .A1(wdata_i[13]),
    .A2(net10));
 sg13g2_a21oi_1 _1633_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1073_),
    .Y(\counter_hi_i.s_count [13]),
    .B1(_1074_));
 sg13g2_inv_1 _1634_ (.VDD(VDD),
    .Y(_1075_),
    .A(_1009_),
    .VSS(VSS));
 sg13g2_nand2_1 _1635_ (.Y(_1076_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .B(_1075_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_2 _1636_ (.VSS(VSS),
    .VDD(VDD),
    .X(_1077_),
    .B(_1076_),
    .A(net27));
 sg13g2_buf_2 fanout59 (.A(net60),
    .X(net59),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1638_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .C(net112),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .Y(_1079_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0972_));
 sg13g2_nor2_1 _1639_ (.A(_1077_),
    .B(_1079_),
    .Y(_1080_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1640_ (.Y(_1081_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .B(_1080_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1641_ (.B1(net7),
    .VDD(VDD),
    .Y(_1082_),
    .VSS(VSS),
    .A1(wdata_i[12]),
    .A2(net10));
 sg13g2_a21oi_1 _1642_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1081_),
    .Y(\counter_hi_i.s_count [12]),
    .B1(_1082_));
 sg13g2_nor2_1 _1643_ (.A(wdata_i[29]),
    .B(net15),
    .Y(_1083_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1644_ (.Y(_1084_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .B(_1015_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1645_ (.Y(_1085_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .B(_1084_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1646_ (.A(net103),
    .B(_1085_),
    .Y(_1086_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1647_ (.A(net74),
    .B(_1083_),
    .C(_1086_),
    .Y(\counter_hi_i.s_count [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1648_ (.B(net112),
    .C(_0972_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .Y(_1087_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1649_ (.A(_1077_),
    .B(_1087_),
    .Y(_1088_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1650_ (.Y(_1089_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .B(_1088_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1651_ (.B1(net9),
    .VDD(VDD),
    .Y(_1090_),
    .VSS(VSS),
    .A1(wdata_i[11]),
    .A2(net12));
 sg13g2_a21oi_1 _1652_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1089_),
    .Y(\counter_hi_i.s_count [11]),
    .B1(_1090_));
 sg13g2_inv_1 _1653_ (.VDD(VDD),
    .Y(_1091_),
    .A(net112),
    .VSS(VSS));
 sg13g2_inv_1 _1654_ (.VDD(VDD),
    .Y(_1092_),
    .A(_0972_),
    .VSS(VSS));
 sg13g2_nor3_1 _1655_ (.A(_1091_),
    .B(_1092_),
    .C(_1077_),
    .Y(_1093_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1656_ (.Y(_1094_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(_1093_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(_0731_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1658_ (.A(wdata_i[10]),
    .B(net18),
    .Y(_1096_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1659_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net14),
    .A2(_1094_),
    .Y(_1097_),
    .B1(_1096_));
 sg13g2_and2_1 _1660_ (.A(net6),
    .B(_1097_),
    .X(\counter_hi_i.s_count [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1661_ (.A(_1092_),
    .B(_1077_),
    .Y(_1098_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1662_ (.Y(_1099_),
    .A(net112),
    .B(_1098_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1663_ (.B1(net9),
    .VDD(VDD),
    .Y(_1100_),
    .VSS(VSS),
    .A1(wdata_i[9]),
    .A2(net12));
 sg13g2_a21oi_1 _1664_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net16),
    .A2(_1099_),
    .Y(\counter_hi_i.s_count [9]),
    .B1(_1100_));
 sg13g2_nor2_1 _1665_ (.A(wdata_i[8]),
    .B(net14),
    .Y(_1101_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1666_ (.Y(_1102_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1667_ (.A(_1102_),
    .B(net27),
    .C(_1076_),
    .Y(_1103_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1668_ (.B(_1103_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .X(_1104_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1669_ (.A(net104),
    .B(_1104_),
    .Y(_1105_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1670_ (.A(net76),
    .B(_1101_),
    .C(_1105_),
    .Y(\counter_hi_i.s_count [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1671_ (.VDD(VDD),
    .Y(_1106_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .VSS(VSS));
 sg13g2_nor2_2 _1672_ (.A(_1106_),
    .B(_1077_),
    .Y(_1107_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1673_ (.B(_1107_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .X(_1108_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1674_ (.A(net104),
    .B(_1108_),
    .Y(_1109_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1675_ (.A(wdata_i[7]),
    .B(_1018_),
    .C(_1019_),
    .Y(_1110_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1676_ (.A(net76),
    .B(_1109_),
    .C(_1110_),
    .Y(\counter_hi_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1677_ (.A(wdata_i[6]),
    .B(net14),
    .Y(_1111_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1678_ (.Y(_1112_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(_1077_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1679_ (.A(net104),
    .B(_1112_),
    .Y(_1113_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1680_ (.A(net75),
    .B(_1111_),
    .C(_1113_),
    .Y(\counter_hi_i.s_count [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1681_ (.A(wdata_i[5]),
    .B(net18),
    .Y(_1114_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 _1682_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .B(net27),
    .C(net106),
    .X(_1115_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1683_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .VDD(VDD),
    .Y(_1116_),
    .VSS(VSS),
    .A1(net27),
    .A2(net106));
 sg13g2_and3_1 _1684_ (.X(_1117_),
    .A(net12),
    .B(_1115_),
    .C(_1116_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1685_ (.A(net75),
    .B(_1114_),
    .C(_1117_),
    .Y(\counter_hi_i.s_count [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1686_ (.A(wdata_i[4]),
    .B(net14),
    .Y(_1118_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 _1687_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .B(net26),
    .C(_1008_),
    .X(_1119_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1688_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .VDD(VDD),
    .Y(_1120_),
    .VSS(VSS),
    .A1(net27),
    .A2(_1008_));
 sg13g2_and3_1 _1689_ (.X(_1121_),
    .A(net11),
    .B(_1119_),
    .C(_1120_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1690_ (.A(net75),
    .B(_1118_),
    .C(_1121_),
    .Y(\counter_hi_i.s_count [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1691_ (.A(wdata_i[3]),
    .B(net18),
    .Y(_1122_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1692_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .C(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .Y(_1123_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 _1693_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .B(net26),
    .C(_1123_),
    .X(_1124_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1694_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .VDD(VDD),
    .Y(_1125_),
    .VSS(VSS),
    .A1(net27),
    .A2(_1123_));
 sg13g2_and3_1 _1695_ (.X(_1126_),
    .A(net11),
    .B(_1124_),
    .C(_1125_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1696_ (.A(net75),
    .B(_1122_),
    .C(_1126_),
    .Y(\counter_hi_i.s_count [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1697_ (.A(wdata_i[2]),
    .B(net18),
    .Y(_1127_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1698_ (.Y(_1128_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 _1699_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(net26),
    .C(_1128_),
    .X(_1129_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1700_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .VDD(VDD),
    .Y(_1130_),
    .VSS(VSS),
    .A1(net26),
    .A2(_1128_));
 sg13g2_and3_1 _1701_ (.X(_1131_),
    .A(net13),
    .B(_1129_),
    .C(_1130_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1702_ (.A(net75),
    .B(_1127_),
    .C(_1131_),
    .Y(\counter_hi_i.s_count [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1703_ (.Y(_1132_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .B(_1015_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1704_ (.B1(net9),
    .VDD(VDD),
    .Y(_1133_),
    .VSS(VSS),
    .A1(wdata_i[28]),
    .A2(net11));
 sg13g2_a21oi_1 _1705_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net15),
    .A2(_1132_),
    .Y(\counter_hi_i.s_count [28]),
    .B1(_1133_));
 sg13g2_nor2_1 _1706_ (.A(wdata_i[1]),
    .B(net18),
    .Y(_1134_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1707_ (.VDD(VDD),
    .Y(_1135_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .VSS(VSS));
 sg13g2_or3_1 _1708_ (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .B(_1135_),
    .C(net26),
    .X(_1136_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1709_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .VDD(VDD),
    .Y(_1137_),
    .VSS(VSS),
    .A1(_1135_),
    .A2(net26));
 sg13g2_and3_1 _1710_ (.X(_1138_),
    .A(net11),
    .B(_1136_),
    .C(_1137_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1711_ (.A(net75),
    .B(_1134_),
    .C(_1138_),
    .Y(\counter_hi_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1712_ (.A(wdata_i[0]),
    .B(net18),
    .Y(_1139_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _1713_ (.A(addr_i[4]),
    .B(addr_i[5]),
    .C(_0937_),
    .Y(_1140_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1714_ (.VDD(VDD),
    .Y(_1141_),
    .A(_1019_),
    .VSS(VSS));
 sg13g2_nor2b_1 _1715_ (.A(net26),
    .B_N(\counter_hi_i.enable_count_i_$_MUX__S_31_B [0]),
    .Y(_1142_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 _1716_ (.VSS(VSS),
    .VDD(VDD),
    .B2(_1141_),
    .C1(_1142_),
    .B1(_1140_),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .Y(_1143_),
    .A2(net26));
 sg13g2_nor3_1 _1717_ (.A(net75),
    .B(_1139_),
    .C(_1143_),
    .Y(\counter_hi_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _1718_ (.A(_0976_),
    .B(net28),
    .C(net106),
    .Y(_1144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1719_ (.Y(_1145_),
    .A(_1144_),
    .B(_1013_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1720_ (.B(_1145_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .X(_1146_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1721_ (.B1(net7),
    .VDD(VDD),
    .Y(_1147_),
    .VSS(VSS),
    .A1(wdata_i[27]),
    .A2(net10));
 sg13g2_a21oi_1 _1722_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net15),
    .A2(_1146_),
    .Y(\counter_hi_i.s_count [27]),
    .B1(_1147_));
 sg13g2_inv_1 _1723_ (.VDD(VDD),
    .Y(_1148_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .VSS(VSS));
 sg13g2_nand3_1 _1724_ (.B(_1144_),
    .C(_1012_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .Y(_1149_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1725_ (.A(_1148_),
    .B(_1149_),
    .Y(_1150_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1726_ (.Y(_1151_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .B(_1150_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1727_ (.Y(_1152_),
    .A(net15),
    .B(_1151_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1728_ (.VDD(VDD),
    .Y(_1153_),
    .A(wdata_i[26]),
    .VSS(VSS));
 sg13g2_a21oi_1 _1729_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1153_),
    .A2(net103),
    .Y(_1154_),
    .B1(net74));
 sg13g2_and2_1 _1730_ (.A(_1152_),
    .B(_1154_),
    .X(\counter_hi_i.s_count [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1731_ (.Y(_1155_),
    .A(_1148_),
    .B(_1149_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1732_ (.B1(net8),
    .VDD(VDD),
    .Y(_1156_),
    .VSS(VSS),
    .A1(wdata_i[25]),
    .A2(net11));
 sg13g2_a21oi_1 _1733_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net15),
    .A2(_1155_),
    .Y(\counter_hi_i.s_count [25]),
    .B1(_1156_));
 sg13g2_nor2_1 _1734_ (.A(wdata_i[24]),
    .B(net15),
    .Y(_1157_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1735_ (.Y(_1158_),
    .A(_1144_),
    .B(_1012_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1736_ (.Y(_1159_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .B(_1158_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1737_ (.A(net103),
    .B(_1159_),
    .Y(_1160_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1738_ (.A(net74),
    .B(_1157_),
    .C(_1160_),
    .Y(\counter_hi_i.s_count [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1739_ (.Y(_1161_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(_1144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1740_ (.B(_1161_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .X(_1162_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1741_ (.B1(net7),
    .VDD(VDD),
    .Y(_1163_),
    .VSS(VSS),
    .A1(wdata_i[23]),
    .A2(net10));
 sg13g2_a21oi_1 _1742_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net15),
    .A2(_1162_),
    .Y(\counter_hi_i.s_count [23]),
    .B1(_1163_));
 sg13g2_xnor2_1 _1743_ (.Y(_1164_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(_1144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1744_ (.Y(_1165_),
    .A(net14),
    .B(_1164_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1745_ (.B1(_1165_),
    .VDD(VDD),
    .Y(_1166_),
    .VSS(VSS),
    .A1(wdata_i[22]),
    .A2(net12));
 sg13g2_nor2_1 _1746_ (.A(net74),
    .B(_1166_),
    .Y(\counter_hi_i.s_count [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1747_ (.B(\counter_hi_i.s_count [30]),
    .A(\counter_hi_i.compare_value_i [30]),
    .X(_1167_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1748_ (.B(\counter_hi_i.s_count [29]),
    .A(\counter_hi_i.compare_value_i [29]),
    .X(_1168_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1749_ (.B(\counter_hi_i.s_count [22]),
    .A(\counter_hi_i.compare_value_i [22]),
    .X(_1169_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1750_ (.B(\counter_hi_i.s_count [10]),
    .A(\counter_hi_i.compare_value_i [10]),
    .X(_1170_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1751_ (.B(\counter_hi_i.s_count [20]),
    .A(\counter_hi_i.compare_value_i [20]),
    .X(_1171_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1752_ (.Y(_1172_),
    .A(net7),
    .B(net10),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(net58),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1754_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .VDD(VDD),
    .Y(_1174_),
    .VSS(VSS),
    .A1(_1018_),
    .A2(_1019_));
 sg13g2_nand3b_1 _1755_ (.B(_1174_),
    .C(net7),
    .Y(_1175_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(_1110_));
 sg13g2_xor2_1 _1756_ (.B(_1175_),
    .A(\counter_hi_i.compare_value_i [7]),
    .X(_1176_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1757_ (.A(net4),
    .B(_1176_),
    .Y(_1177_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1758_ (.A0(_1177_),
    .A1(_1176_),
    .S(_1107_),
    .X(_1178_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _1759_ (.Y(_1179_),
    .B1(_1178_),
    .B2(_1088_),
    .A2(_1176_),
    .A1(net4),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1760_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .A2(net18),
    .Y(_1180_),
    .B1(_1090_));
 sg13g2_xnor2_1 _1761_ (.Y(_1181_),
    .A(\counter_hi_i.compare_value_i [11]),
    .B(_1180_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _1762_ (.A(_1179_),
    .B_N(_1181_),
    .Y(_1182_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1763_ (.B(_1176_),
    .A(_1107_),
    .X(_1183_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1764_ (.A(_1088_),
    .B(net4),
    .C(_1181_),
    .D(_1183_),
    .Y(_1184_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1765_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .A2(net13),
    .Y(_1185_),
    .B1(_1051_));
 sg13g2_xor2_1 _1766_ (.B(_1185_),
    .A(\counter_hi_i.compare_value_i [19]),
    .X(_1186_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1767_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .VDD(VDD),
    .Y(_1187_),
    .VSS(VSS),
    .A1(_1018_),
    .A2(_1019_));
 sg13g2_nand3b_1 _1768_ (.B(_1187_),
    .C(net7),
    .Y(_1188_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(_1041_));
 sg13g2_xor2_1 _1769_ (.B(_1188_),
    .A(\counter_hi_i.compare_value_i [21]),
    .X(_1189_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1770_ (.A(net3),
    .B(_1189_),
    .Y(_1190_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1771_ (.A0(_1189_),
    .A1(_1190_),
    .S(_0964_),
    .X(_1191_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _1772_ (.Y(_1192_),
    .B1(_1191_),
    .B2(_1047_),
    .A2(_1189_),
    .A1(net4),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _1773_ (.B(_1186_),
    .C(_1190_),
    .Y(_1193_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(_1047_));
 sg13g2_o21ai_1 _1774_ (.B1(_1193_),
    .VDD(VDD),
    .Y(_1194_),
    .VSS(VSS),
    .A1(_1186_),
    .A2(_1192_));
 sg13g2_o21ai_1 _1775_ (.B1(_1194_),
    .VDD(VDD),
    .Y(_1195_),
    .VSS(VSS),
    .A1(_1182_),
    .A2(_1184_));
 sg13g2_or4_1 _1776_ (.A(_1169_),
    .B(_1170_),
    .C(_1171_),
    .D(_1195_),
    .X(_1196_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1777_ (.Y(_1197_),
    .A(\counter_hi_i.compare_value_i [31]),
    .B(\counter_hi_i.s_count [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1778_ (.B(\counter_hi_i.s_count [6]),
    .A(\counter_hi_i.compare_value_i [6]),
    .X(_1198_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1779_ (.A(_1063_),
    .B(_0974_),
    .Y(_1199_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1780_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .A2(net13),
    .Y(_1200_),
    .B1(_1082_));
 sg13g2_xnor2_1 _1781_ (.Y(_1201_),
    .A(\counter_hi_i.compare_value_i [12]),
    .B(_1200_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1782_ (.B1(_1201_),
    .VDD(VDD),
    .Y(_1202_),
    .VSS(VSS),
    .A1(net3),
    .A2(_1199_));
 sg13g2_a21oi_1 _1783_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .A2(net17),
    .Y(_1203_),
    .B1(_1069_));
 sg13g2_xnor2_1 _1784_ (.Y(_1204_),
    .A(\counter_hi_i.compare_value_i [15]),
    .B(_1203_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1785_ (.Y(_1205_),
    .A(_1202_),
    .B(_1204_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1786_ (.Y(_1206_),
    .A(\counter_hi_i.compare_value_i [14]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1787_ (.VDD(VDD),
    .Y(_1207_),
    .A(_1206_),
    .VSS(VSS));
 sg13g2_nor3_1 _1788_ (.A(_1070_),
    .B(net3),
    .C(_1207_),
    .Y(_1208_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1789_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .C(_1064_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .Y(_1209_),
    .VDD(VDD),
    .VSS(VSS),
    .D(net12));
 sg13g2_nor2b_1 _1790_ (.A(_1072_),
    .B_N(_1209_),
    .Y(_1210_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1791_ (.B(_1064_),
    .C(net10),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .Y(_1211_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1792_ (.Y(_1212_),
    .A(wdata_i[14]),
    .B(net104),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1793_ (.B1(_1212_),
    .VDD(VDD),
    .Y(_1213_),
    .VSS(VSS),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .A2(_1211_));
 sg13g2_nand3_1 _1794_ (.B(net6),
    .C(_1213_),
    .A(\counter_hi_i.compare_value_i [14]),
    .Y(_1214_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1795_ (.B1(_1214_),
    .VDD(VDD),
    .Y(_0122_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [14]),
    .A2(_1210_));
 sg13g2_nor2_1 _1796_ (.A(_1208_),
    .B(_0122_),
    .Y(_0123_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _1797_ (.A(net74),
    .B(net104),
    .Y(_0124_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1798_ (.Y(_0125_),
    .A(_0124_),
    .B(_1207_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1799_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .A2(net13),
    .Y(_0126_),
    .B1(_1163_));
 sg13g2_xnor2_1 _1800_ (.Y(_0127_),
    .A(\counter_hi_i.compare_value_i [23]),
    .B(_0126_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1801_ (.B(_0124_),
    .C(_0127_),
    .A(_1161_),
    .Y(_0128_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1802_ (.B1(_0128_),
    .VDD(VDD),
    .Y(_0129_),
    .VSS(VSS),
    .A1(_1065_),
    .A2(_0125_));
 sg13g2_nand3_1 _1803_ (.B(wdata_i[22]),
    .C(net6),
    .A(\counter_hi_i.compare_value_i [22]),
    .Y(_0130_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1804_ (.B1(_0130_),
    .VDD(VDD),
    .Y(_0131_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [22]),
    .A2(wdata_i[22]));
 sg13g2_nand3_1 _1805_ (.B(_1013_),
    .C(net10),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .Y(_0132_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1806_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net8),
    .A2(_0132_),
    .Y(_0133_),
    .B1(\counter_hi_i.compare_value_i [22]));
 sg13g2_a21oi_1 _1807_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net103),
    .A2(_0131_),
    .Y(_0134_),
    .B1(_0133_));
 sg13g2_a21oi_1 _1808_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .A2(net13),
    .Y(_0135_),
    .B1(_1147_));
 sg13g2_xor2_1 _1809_ (.B(_0135_),
    .A(\counter_hi_i.compare_value_i [27]),
    .X(_0136_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1810_ (.Y(_0137_),
    .A(_0134_),
    .B(_0136_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1811_ (.B1(_0137_),
    .VDD(VDD),
    .Y(_0138_),
    .VSS(VSS),
    .A1(_1161_),
    .A2(_0127_));
 sg13g2_or4_1 _1812_ (.A(_1205_),
    .B(_0123_),
    .C(_0129_),
    .D(_0138_),
    .X(_0139_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1813_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .A2(net17),
    .Y(_0140_),
    .B1(_1053_));
 sg13g2_xnor2_1 _1814_ (.Y(_0141_),
    .A(\counter_hi_i.compare_value_i [18]),
    .B(_0140_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1815_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .A(\counter_hi_i.compare_value_i [17]),
    .X(_0142_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1816_ (.A(net3),
    .B(_0142_),
    .Y(_0143_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1817_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .A2(net13),
    .Y(_0144_),
    .B1(_1074_));
 sg13g2_xnor2_1 _1818_ (.Y(_0145_),
    .A(\counter_hi_i.compare_value_i [13]),
    .B(_0144_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1819_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1066_),
    .A2(_0143_),
    .Y(_0146_),
    .B1(_0145_));
 sg13g2_or2_1 _1820_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0147_),
    .B(_0146_),
    .A(_0141_));
 sg13g2_o21ai_1 _1821_ (.B1(_0145_),
    .VDD(VDD),
    .Y(_0148_),
    .VSS(VSS),
    .A1(_1038_),
    .A2(net4));
 sg13g2_a21oi_1 _1822_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .A2(net17),
    .Y(_0149_),
    .B1(_1058_));
 sg13g2_xnor2_1 _1823_ (.Y(_0150_),
    .A(\counter_hi_i.compare_value_i [17]),
    .B(_0149_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1824_ (.A0(_0143_),
    .A1(_0150_),
    .S(_0969_),
    .X(_0151_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1825_ (.A(\counter_hi_i.compare_value_i [17]),
    .B(wdata_i[17]),
    .Y(_0152_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _1826_ (.X(_0153_),
    .A(\counter_hi_i.compare_value_i [17]),
    .B(wdata_i[17]),
    .C(net8),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1827_ (.B1(net103),
    .VDD(VDD),
    .Y(_0154_),
    .VSS(VSS),
    .A1(_0152_),
    .A2(_0153_));
 sg13g2_nand2b_1 _1828_ (.Y(_0155_),
    .B(net74),
    .A_N(\counter_hi_i.compare_value_i [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1829_ (.B(_0154_),
    .C(_0155_),
    .A(_0145_),
    .Y(_0156_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1830_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1055_),
    .A2(_0151_),
    .Y(_0157_),
    .B1(_0156_));
 sg13g2_a21o_1 _1831_ (.A2(_0148_),
    .A1(_0147_),
    .B1(_0157_),
    .X(_0158_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1832_ (.Y(_0159_),
    .A(\counter_hi_i.compare_value_i [25]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1833_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .A(\counter_hi_i.compare_value_i [26]),
    .X(_0160_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1834_ (.A(net3),
    .B(_0160_),
    .Y(_0161_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1835_ (.B(_0159_),
    .C(_0161_),
    .A(_1149_),
    .Y(_0162_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1836_ (.Y(_0163_),
    .A(_1153_),
    .B(net103),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1837_ (.Y(_0164_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .B(net10),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _1838_ (.A(\counter_hi_i.compare_value_i [26]),
    .B(net8),
    .C(_0163_),
    .D(_0164_),
    .X(_0165_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1839_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1154_),
    .A2(_0164_),
    .Y(_0166_),
    .B1(\counter_hi_i.compare_value_i [26]));
 sg13g2_o21ai_1 _1840_ (.B1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .Y(_0167_),
    .VSS(VSS),
    .A1(_0165_),
    .A2(_0166_));
 sg13g2_nand2_1 _1841_ (.Y(_0168_),
    .A(_1148_),
    .B(_0161_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1842_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_0167_),
    .A2(_0168_),
    .Y(_0169_),
    .B1(_1149_));
 sg13g2_nand3_1 _1843_ (.B(wdata_i[26]),
    .C(net7),
    .A(\counter_hi_i.compare_value_i [26]),
    .Y(_0170_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1844_ (.B1(_0170_),
    .VDD(VDD),
    .Y(_0171_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [26]),
    .A2(wdata_i[26]));
 sg13g2_nand2_1 _1845_ (.Y(_0172_),
    .A(net103),
    .B(_0171_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1846_ (.B1(_0172_),
    .VDD(VDD),
    .Y(_0173_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [26]),
    .A2(net6));
 sg13g2_a21oi_1 _1847_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .A2(net18),
    .Y(_0174_),
    .B1(_1156_));
 sg13g2_xnor2_1 _1848_ (.Y(_0175_),
    .A(\counter_hi_i.compare_value_i [25]),
    .B(_0174_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1849_ (.B1(_0175_),
    .VDD(VDD),
    .Y(_0176_),
    .VSS(VSS),
    .A1(_0169_),
    .A2(_0173_));
 sg13g2_xor2_1 _1850_ (.B(\counter_hi_i.s_count [2]),
    .A(\counter_hi_i.compare_value_i [2]),
    .X(_0177_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _1851_ (.A2(_0176_),
    .A1(_0162_),
    .B1(_0177_),
    .X(_0178_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1852_ (.A(_1198_),
    .B(_0139_),
    .C(_0158_),
    .D(_0178_),
    .Y(_0179_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1853_ (.B(wdata_i[9]),
    .C(net6),
    .A(\counter_hi_i.compare_value_i [9]),
    .Y(_0180_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1854_ (.B1(_0180_),
    .VDD(VDD),
    .Y(_0181_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [9]),
    .A2(wdata_i[9]));
 sg13g2_nand2_1 _1855_ (.Y(_0182_),
    .A(net104),
    .B(_0181_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1856_ (.B1(_0182_),
    .VDD(VDD),
    .Y(_0183_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [9]),
    .A2(net6));
 sg13g2_xor2_1 _1857_ (.B(net112),
    .A(\counter_hi_i.compare_value_i [9]),
    .X(_0184_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1858_ (.A(net3),
    .B(_0184_),
    .Y(_0185_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1859_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net112),
    .A2(net17),
    .Y(_0186_),
    .B1(_1100_));
 sg13g2_nor2_1 _1860_ (.A(wdata_i[9]),
    .B(net17),
    .Y(_0187_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1861_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net112),
    .A2(net13),
    .Y(_0188_),
    .B1(_0187_));
 sg13g2_nand3_1 _1862_ (.B(net6),
    .C(_0188_),
    .A(\counter_hi_i.compare_value_i [9]),
    .Y(_0189_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1863_ (.B1(_0189_),
    .VDD(VDD),
    .Y(_0190_),
    .VSS(VSS),
    .A1(\counter_hi_i.compare_value_i [9]),
    .A2(_0186_));
 sg13g2_mux2_1 _1864_ (.A0(_0185_),
    .A1(_0190_),
    .S(_0972_),
    .X(_0191_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _1865_ (.Y(_0192_),
    .B(_1201_),
    .A_N(_1079_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1866_ (.Y(_0193_),
    .A(\counter_hi_i.compare_value_i [12]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1867_ (.B(_1079_),
    .C(_0124_),
    .A(_0972_),
    .Y(_0194_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0193_));
 sg13g2_a21oi_1 _1868_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_0192_),
    .A2(_0194_),
    .Y(_0195_),
    .B1(_1077_));
 sg13g2_nand2_1 _1869_ (.Y(_0196_),
    .A(_0193_),
    .B(_0185_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1870_ (.A(_1098_),
    .B(_0196_),
    .Y(_0197_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 _1871_ (.VSS(VSS),
    .VDD(VDD),
    .B2(_0195_),
    .C1(_0197_),
    .B1(_0191_),
    .A1(_1201_),
    .Y(_0198_),
    .A2(_0183_));
 sg13g2_xor2_1 _1872_ (.B(\counter_hi_i.s_count [8]),
    .A(\counter_hi_i.compare_value_i [8]),
    .X(_0199_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1873_ (.A(\counter_hi_i.compare_value_i [24]),
    .B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .C(net74),
    .Y(_0200_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1874_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.compare_value_i [24]),
    .A2(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .Y(_0201_),
    .B1(_0200_));
 sg13g2_nand2_1 _1875_ (.Y(_0202_),
    .A(_1012_),
    .B(net12),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1876_ (.A(_0976_),
    .B(_0201_),
    .C(_0202_),
    .Y(_0203_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1877_ (.A(_0970_),
    .B(_0975_),
    .C(_0141_),
    .Y(_0204_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1878_ (.B1(_1065_),
    .VDD(VDD),
    .Y(_0205_),
    .VSS(VSS),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_xor2_1 _1879_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .A(\counter_hi_i.compare_value_i [24]),
    .X(_0206_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1880_ (.B(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .C(_1144_),
    .A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .Y(_0207_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1881_ (.B(_0206_),
    .C(_0207_),
    .A(_0124_),
    .Y(_0208_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1882_ (.Y(_0209_),
    .A(\counter_hi_i.compare_value_i [0]),
    .B(\counter_hi_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1883_ (.Y(_0210_),
    .A(wdata_i[24]),
    .B(net6),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1884_ (.B(_0210_),
    .A(\counter_hi_i.compare_value_i [24]),
    .X(_0211_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1885_ (.B(_0127_),
    .C(_0211_),
    .A(_0141_),
    .Y(_0212_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1886_ (.A(_0976_),
    .B(_1014_),
    .Y(_0213_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1887_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_1065_),
    .A2(_0213_),
    .Y(_0214_),
    .B1(net3));
 sg13g2_a21oi_1 _1888_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .A2(net13),
    .Y(_0215_),
    .B1(_1133_));
 sg13g2_xnor2_1 _1889_ (.Y(_0216_),
    .A(\counter_hi_i.compare_value_i [28]),
    .B(_0215_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1890_ (.Y(_0217_),
    .A(_0214_),
    .B(_0216_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1891_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net3),
    .A2(_0212_),
    .Y(_0218_),
    .B1(_0217_));
 sg13g2_nand4_1 _1892_ (.B(_0208_),
    .C(_0209_),
    .A(_0205_),
    .Y(_0219_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0218_));
 sg13g2_nor3_1 _1893_ (.A(_0198_),
    .B(_0199_),
    .C(_0219_),
    .Y(_0220_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1894_ (.Y(_0221_),
    .A(\counter_hi_i.compare_value_i [16]),
    .B(\counter_hi_i.s_count [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1895_ (.B(\counter_hi_i.s_count [4]),
    .A(\counter_hi_i.compare_value_i [4]),
    .X(_0222_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1896_ (.B(\counter_hi_i.s_count [1]),
    .A(\counter_hi_i.compare_value_i [1]),
    .X(_0223_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1897_ (.B(\counter_hi_i.s_count [3]),
    .A(\counter_hi_i.compare_value_i [3]),
    .X(_0224_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1898_ (.B(\counter_hi_i.s_count [5]),
    .A(\counter_hi_i.compare_value_i [5]),
    .X(_0225_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _1899_ (.A(_0222_),
    .B(_0223_),
    .C(_0224_),
    .D(_0225_),
    .Y(_0226_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _1900_ (.A(_0221_),
    .B(_0226_),
    .X(_0227_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1901_ (.B(_0179_),
    .C(_0220_),
    .A(_1197_),
    .Y(_0228_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0227_));
 sg13g2_nor4_1 _1902_ (.A(_1167_),
    .B(_1168_),
    .C(_1196_),
    .D(_0228_),
    .Y(\counter_hi_i.target_reached_o_reg_D ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _1903_ (.A(addr_i[2]),
    .B(addr_i[3]),
    .C(addr_i[0]),
    .Y(_0229_),
    .VDD(VDD),
    .VSS(VSS),
    .D(addr_i[1]));
 sg13g2_nand2_2 _1904_ (.Y(_0230_),
    .A(_0938_),
    .B(_0229_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1906_ (.A0(wdata_i[0]),
    .A1(\counter_lo_i.compare_value_i [0]),
    .S(net101),
    .X(_0032_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1907_ (.A0(wdata_i[10]),
    .A1(\counter_lo_i.compare_value_i [10]),
    .S(net102),
    .X(_0033_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1908_ (.A0(wdata_i[11]),
    .A1(\counter_lo_i.compare_value_i [11]),
    .S(net102),
    .X(_0034_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1909_ (.A0(wdata_i[12]),
    .A1(\counter_lo_i.compare_value_i [12]),
    .S(net102),
    .X(_0035_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1910_ (.A0(wdata_i[13]),
    .A1(\counter_lo_i.compare_value_i [13]),
    .S(net102),
    .X(_0036_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1911_ (.A0(wdata_i[14]),
    .A1(\counter_lo_i.compare_value_i [14]),
    .S(net99),
    .X(_0037_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout55 (.A(net58),
    .X(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1913_ (.A0(wdata_i[15]),
    .A1(\counter_lo_i.compare_value_i [15]),
    .S(net100),
    .X(_0038_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1914_ (.A0(wdata_i[16]),
    .A1(\counter_lo_i.compare_value_i [16]),
    .S(net100),
    .X(_0039_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1915_ (.A0(wdata_i[17]),
    .A1(\counter_lo_i.compare_value_i [17]),
    .S(net99),
    .X(_0040_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1916_ (.A0(wdata_i[18]),
    .A1(\counter_lo_i.compare_value_i [18]),
    .S(net99),
    .X(_0041_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1917_ (.A0(wdata_i[19]),
    .A1(\counter_lo_i.compare_value_i [19]),
    .S(net99),
    .X(_0042_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1918_ (.VDD(VDD),
    .Y(_0233_),
    .A(wdata_i[1]),
    .VSS(VSS));
 sg13g2_nand2_1 _1919_ (.Y(_0234_),
    .A(\counter_lo_i.compare_value_i [1]),
    .B(net101),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1920_ (.B1(_0234_),
    .VDD(VDD),
    .Y(_0043_),
    .VSS(VSS),
    .A1(_0233_),
    .A2(net101));
 sg13g2_mux2_1 _1921_ (.A0(wdata_i[20]),
    .A1(\counter_lo_i.compare_value_i [20]),
    .S(net99),
    .X(_0044_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1922_ (.A0(wdata_i[21]),
    .A1(\counter_lo_i.compare_value_i [21]),
    .S(net98),
    .X(_0045_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1923_ (.A0(wdata_i[22]),
    .A1(\counter_lo_i.compare_value_i [22]),
    .S(net98),
    .X(_0046_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1924_ (.A0(wdata_i[23]),
    .A1(\counter_lo_i.compare_value_i [23]),
    .S(net98),
    .X(_0047_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1925_ (.A0(wdata_i[24]),
    .A1(\counter_lo_i.compare_value_i [24]),
    .S(net99),
    .X(_0048_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(net58),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1927_ (.A0(wdata_i[25]),
    .A1(\counter_lo_i.compare_value_i [25]),
    .S(net98),
    .X(_0049_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1928_ (.Y(_0236_),
    .A(\counter_lo_i.compare_value_i [26]),
    .B(net99),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _1929_ (.B1(_0236_),
    .VDD(VDD),
    .Y(_0050_),
    .VSS(VSS),
    .A1(_1153_),
    .A2(net99));
 sg13g2_mux2_1 _1930_ (.A0(wdata_i[27]),
    .A1(\counter_lo_i.compare_value_i [27]),
    .S(net100),
    .X(_0051_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1931_ (.A0(wdata_i[28]),
    .A1(\counter_lo_i.compare_value_i [28]),
    .S(net98),
    .X(_0052_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1932_ (.A0(wdata_i[29]),
    .A1(\counter_lo_i.compare_value_i [29]),
    .S(net98),
    .X(_0053_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1933_ (.A0(wdata_i[2]),
    .A1(\counter_lo_i.compare_value_i [2]),
    .S(net101),
    .X(_0054_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1934_ (.A0(wdata_i[30]),
    .A1(\counter_lo_i.compare_value_i [30]),
    .S(net98),
    .X(_0055_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1935_ (.A0(wdata_i[31]),
    .A1(\counter_lo_i.compare_value_i [31]),
    .S(net98),
    .X(_0056_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1936_ (.A0(wdata_i[3]),
    .A1(\counter_lo_i.compare_value_i [3]),
    .S(net101),
    .X(_0057_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1937_ (.A0(wdata_i[4]),
    .A1(\counter_lo_i.compare_value_i [4]),
    .S(net101),
    .X(_0058_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1938_ (.A0(wdata_i[5]),
    .A1(\counter_lo_i.compare_value_i [5]),
    .S(net101),
    .X(_0059_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1939_ (.A0(wdata_i[6]),
    .A1(\counter_lo_i.compare_value_i [6]),
    .S(net101),
    .X(_0060_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1940_ (.A0(wdata_i[7]),
    .A1(\counter_lo_i.compare_value_i [7]),
    .S(net102),
    .X(_0061_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1941_ (.A0(wdata_i[8]),
    .A1(\counter_lo_i.compare_value_i [8]),
    .S(net102),
    .X(_0062_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _1942_ (.A0(wdata_i[9]),
    .A1(\counter_lo_i.compare_value_i [9]),
    .S(net102),
    .X(_0063_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1943_ (.VDD(VDD),
    .Y(_0237_),
    .A(s_cfg_lo_reg[4]),
    .VSS(VSS));
 sg13g2_inv_1 _1944_ (.VDD(VDD),
    .Y(_0238_),
    .A(s_cfg_lo_reg[31]),
    .VSS(VSS));
 sg13g2_o21ai_1 _1945_ (.B1(\counter_lo_i.target_reached_o ),
    .VDD(VDD),
    .Y(_0239_),
    .VSS(VSS),
    .A1(_0238_),
    .A2(\counter_hi_i.target_reached_o ));
 sg13g2_and2_1 _1946_ (.A(_0957_),
    .B(_0958_),
    .X(_0240_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_2 _1947_ (.VSS(VSS),
    .VDD(VDD),
    .B1(s_cfg_lo_reg[1]),
    .Y(_0241_),
    .A2(_0229_),
    .A1(_0240_));
 sg13g2_o21ai_1 _1948_ (.B1(_0241_),
    .VDD(VDD),
    .Y(_0242_),
    .VSS(VSS),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(_0734_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(net53),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _1951_ (.Y(_0245_),
    .A(addr_i[3]),
    .B(_0939_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1952_ (.A(addr_i[2]),
    .B(_0245_),
    .Y(_0246_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 _1953_ (.Y(_0247_),
    .A(_1140_),
    .B(_0246_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(net52),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(net53),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1956_ (.A(wdata_i[31]),
    .B(net66),
    .Y(_0250_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1957_ (.VDD(VDD),
    .Y(_0251_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .VSS(VSS));
 sg13g2_inv_1 _1958_ (.VDD(VDD),
    .Y(_0252_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .VSS(VSS));
 sg13g2_nand3_1 _1959_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .C(\counter_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .Y(_0253_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1960_ (.A(_0252_),
    .B(_0253_),
    .Y(_0254_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1961_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .C(_0254_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .Y(_0255_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _1962_ (.X(_0256_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .C(\counter_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _1963_ (.X(_0257_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .C(_0256_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1964_ (.VDD(VDD),
    .Y(_0258_),
    .A(\counter_lo_i.enable_count_i_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_B ),
    .VSS(VSS));
 sg13g2_nand4_1 _1965_ (.B(_0258_),
    .C(s_cfg_lo_reg[7]),
    .A(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ),
    .Y(_0259_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0978_));
 sg13g2_and4_1 _1966_ (.A(\counter_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .C(_1000_),
    .D(_0259_),
    .X(_0260_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(net53),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _1968_ (.A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .C(\counter_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .D(\counter_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .X(_0262_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _1969_ (.B(_0257_),
    .C(net5),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .Y(_0263_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0262_));
 sg13g2_buf_2 fanout48 (.A(_0737_),
    .X(net48),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _1971_ (.VDD(VDD),
    .Y(_0265_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .VSS(VSS));
 sg13g2_nand2_1 _1972_ (.Y(_0266_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1973_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .C(\counter_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .Y(_0267_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1974_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .C(\counter_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .Y(_0268_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _1975_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0269_),
    .B(_0268_),
    .A(_0267_));
 sg13g2_nor3_2 _1976_ (.A(_0265_),
    .B(_0266_),
    .C(_0269_),
    .Y(_0270_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1977_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .C(_0270_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .Y(_0271_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _1978_ (.A(_0251_),
    .B(_0255_),
    .C(net19),
    .Y(_0272_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0271_));
 sg13g2_nand2_1 _1979_ (.Y(_0273_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .B(_0272_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1980_ (.Y(_0274_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [31]),
    .B(_0273_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1981_ (.A(addr_i[2]),
    .B(_1018_),
    .C(_0245_),
    .Y(_0275_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout46 (.A(net48),
    .X(net46),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1984_ (.A(_0274_),
    .B(net94),
    .Y(_0278_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1985_ (.A(net71),
    .B(_0250_),
    .C(_0278_),
    .Y(\counter_lo_i.s_count [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1986_ (.A(wdata_i[30]),
    .B(net64),
    .Y(_0279_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _1987_ (.B(_0272_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .X(_0280_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1988_ (.A(net94),
    .B(_0280_),
    .Y(_0281_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _1989_ (.A(net69),
    .B(_0279_),
    .C(_0281_),
    .Y(\counter_lo_i.s_count [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout45 (.A(net48),
    .X(net45),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout44 (.A(net48),
    .X(net44),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _1992_ (.A(_0255_),
    .B(net19),
    .C(_0267_),
    .Y(_0284_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _1993_ (.Y(_0285_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .B(_0284_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1994_ (.A(wdata_i[21]),
    .B(net64),
    .Y(_0286_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _1995_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net64),
    .A2(_0285_),
    .Y(_0287_),
    .B1(_0286_));
 sg13g2_nor2b_1 _1996_ (.A(net69),
    .B_N(_0287_),
    .Y(\counter_lo_i.s_count [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1997_ (.A(wdata_i[20]),
    .B(net65),
    .Y(_0288_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _1998_ (.A(_0255_),
    .B(net20),
    .Y(_0289_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _1999_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .C(_0289_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .Y(_0290_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2000_ (.Y(_0291_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(_0290_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2001_ (.A(net93),
    .B(_0291_),
    .Y(_0292_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2002_ (.A(net70),
    .B(_0288_),
    .C(_0292_),
    .Y(\counter_lo_i.s_count [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2003_ (.A(wdata_i[19]),
    .B(net65),
    .Y(_0293_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2004_ (.VDD(VDD),
    .Y(_0294_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .VSS(VSS));
 sg13g2_nor3_1 _2005_ (.A(_0294_),
    .B(_0255_),
    .C(net19),
    .Y(_0295_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2006_ (.B(_0295_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .X(_0296_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2007_ (.A(net93),
    .B(_0296_),
    .Y(_0297_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2008_ (.A(net70),
    .B(_0293_),
    .C(_0297_),
    .Y(\counter_lo_i.s_count [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2009_ (.A(wdata_i[18]),
    .B(net65),
    .Y(_0298_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout43 (.A(_0739_),
    .X(net43),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2011_ (.Y(_0300_),
    .A(_0294_),
    .B(_0289_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2012_ (.A(net93),
    .B(_0300_),
    .Y(_0301_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2013_ (.A(net70),
    .B(_0298_),
    .C(_0301_),
    .Y(\counter_lo_i.s_count [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2014_ (.A(wdata_i[17]),
    .B(net65),
    .Y(_0302_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2015_ (.Y(_0303_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .B(_0254_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2016_ (.A(_0303_),
    .B(net19),
    .Y(_0304_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2017_ (.B(_0304_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .X(_0305_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2018_ (.A(net93),
    .B(_0305_),
    .Y(_0306_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2019_ (.A(net70),
    .B(_0302_),
    .C(_0306_),
    .Y(\counter_lo_i.s_count [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2020_ (.A(wdata_i[16]),
    .B(net65),
    .Y(_0307_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2021_ (.A(_0252_),
    .B(_0253_),
    .C(net20),
    .Y(_0308_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2022_ (.B(_0308_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .X(_0309_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2023_ (.A(net97),
    .B(_0309_),
    .Y(_0310_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2024_ (.A(net70),
    .B(_0307_),
    .C(_0310_),
    .Y(\counter_lo_i.s_count [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2025_ (.A(wdata_i[15]),
    .B(net65),
    .Y(_0311_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2026_ (.A(_0253_),
    .B(net20),
    .Y(_0312_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2027_ (.Y(_0313_),
    .A(_0252_),
    .B(_0312_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2028_ (.A(net97),
    .B(_0313_),
    .Y(_0314_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2029_ (.A(net70),
    .B(_0311_),
    .C(_0314_),
    .Y(\counter_lo_i.s_count [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2030_ (.A(wdata_i[14]),
    .B(net66),
    .Y(_0315_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2031_ (.VDD(VDD),
    .Y(_0316_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .VSS(VSS));
 sg13g2_inv_1 _2032_ (.VDD(VDD),
    .Y(_0317_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .VSS(VSS));
 sg13g2_nor3_1 _2033_ (.A(_0316_),
    .B(_0317_),
    .C(net20),
    .Y(_0318_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2034_ (.B(_0318_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .X(_0319_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2035_ (.A(net93),
    .B(_0319_),
    .Y(_0320_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2036_ (.A(net71),
    .B(_0315_),
    .C(_0320_),
    .Y(\counter_lo_i.s_count [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2037_ (.A(wdata_i[13]),
    .B(net66),
    .Y(_0321_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2038_ (.A(_0316_),
    .B(net20),
    .Y(_0322_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2039_ (.Y(_0323_),
    .A(_0317_),
    .B(_0322_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2040_ (.A(net93),
    .B(_0323_),
    .Y(_0324_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2041_ (.A(net71),
    .B(_0321_),
    .C(_0324_),
    .Y(\counter_lo_i.s_count [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2042_ (.A(wdata_i[12]),
    .B(net68),
    .Y(_0325_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2043_ (.Y(_0326_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .B(net20),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2044_ (.A(net96),
    .B(_0326_),
    .Y(_0327_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2045_ (.A(_0242_),
    .B(_0325_),
    .C(_0327_),
    .Y(\counter_lo_i.s_count [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2046_ (.A(wdata_i[29]),
    .B(net64),
    .Y(_0328_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2047_ (.A(_0255_),
    .B(net19),
    .C(_0271_),
    .Y(_0329_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2048_ (.Y(_0330_),
    .A(_0251_),
    .B(_0329_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2049_ (.A(net94),
    .B(_0330_),
    .Y(_0331_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2050_ (.A(net69),
    .B(_0328_),
    .C(_0331_),
    .Y(\counter_lo_i.s_count [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2051_ (.A(wdata_i[11]),
    .B(net68),
    .Y(_0332_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2052_ (.VDD(VDD),
    .Y(_0333_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .VSS(VSS));
 sg13g2_inv_1 _2053_ (.VDD(VDD),
    .Y(_0334_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .VSS(VSS));
 sg13g2_nand4_1 _2054_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .C(_0257_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .Y(_0335_),
    .VDD(VDD),
    .VSS(VSS),
    .D(net5));
 sg13g2_nor3_1 _2055_ (.A(_0333_),
    .B(_0334_),
    .C(_0335_),
    .Y(_0336_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2056_ (.B(_0336_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .X(_0337_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2057_ (.A(net96),
    .B(_0337_),
    .Y(_0338_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2058_ (.A(net73),
    .B(_0332_),
    .C(_0338_),
    .Y(\counter_lo_i.s_count [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2059_ (.A(wdata_i[10]),
    .B(net68),
    .Y(_0339_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2060_ (.A(_0334_),
    .B(_0335_),
    .Y(_0340_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2061_ (.Y(_0341_),
    .A(_0333_),
    .B(_0340_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2062_ (.A(net96),
    .B(_0341_),
    .Y(_0342_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2063_ (.A(net73),
    .B(_0339_),
    .C(_0342_),
    .Y(\counter_lo_i.s_count [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2064_ (.Y(_0343_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .B(_0335_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _2065_ (.Y(_0344_),
    .B(net95),
    .A_N(wdata_i[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2066_ (.B1(_0344_),
    .VDD(VDD),
    .Y(_0345_),
    .VSS(VSS),
    .A1(net95),
    .A2(_0343_));
 sg13g2_nor2_1 _2067_ (.A(net73),
    .B(_0345_),
    .Y(\counter_lo_i.s_count [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2068_ (.A(wdata_i[8]),
    .B(net68),
    .Y(_0346_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2069_ (.A(_0257_),
    .B(net5),
    .X(_0347_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2070_ (.Y(_0348_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .B(_0347_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2071_ (.Y(_0349_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(_0348_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2072_ (.A(net96),
    .B(_0349_),
    .Y(_0350_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2073_ (.A(net73),
    .B(_0346_),
    .C(_0350_),
    .Y(\counter_lo_i.s_count [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2074_ (.A(wdata_i[7]),
    .B(net68),
    .Y(_0351_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2075_ (.B(_0347_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .X(_0352_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2076_ (.A(net96),
    .B(_0352_),
    .Y(_0353_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2077_ (.A(net73),
    .B(_0351_),
    .C(_0353_),
    .Y(\counter_lo_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2078_ (.A(wdata_i[6]),
    .B(net67),
    .Y(_0354_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2079_ (.B(_0256_),
    .C(net5),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .Y(_0355_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2080_ (.Y(_0356_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(_0355_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2081_ (.A(net95),
    .B(_0356_),
    .Y(_0357_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2082_ (.A(net72),
    .B(_0354_),
    .C(_0357_),
    .Y(\counter_lo_i.s_count [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2083_ (.A(wdata_i[5]),
    .B(net67),
    .Y(_0358_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2084_ (.Y(_0359_),
    .A(_0256_),
    .B(net5),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2085_ (.Y(_0360_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .B(_0359_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2086_ (.A(net95),
    .B(_0360_),
    .Y(_0361_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2087_ (.A(net72),
    .B(_0358_),
    .C(_0361_),
    .Y(\counter_lo_i.s_count [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2088_ (.A(wdata_i[4]),
    .B(net67),
    .Y(_0362_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2089_ (.B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .C(net5),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .Y(_0363_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2090_ (.Y(_0364_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .B(_0363_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2091_ (.A(net95),
    .B(_0364_),
    .Y(_0365_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2092_ (.A(net72),
    .B(_0362_),
    .C(_0365_),
    .Y(\counter_lo_i.s_count [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _2093_ (.Y(_0366_),
    .B(net95),
    .A_N(wdata_i[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2094_ (.VDD(VDD),
    .Y(_0367_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .VSS(VSS));
 sg13g2_nand3_1 _2095_ (.B(_0367_),
    .C(net5),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .Y(_0368_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _2096_ (.A2(_0260_),
    .A1(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .B1(_0367_),
    .X(_0369_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2097_ (.B(_0368_),
    .C(_0369_),
    .A(net67),
    .Y(_0370_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2098_ (.A(_0366_),
    .B(_0370_),
    .X(_0371_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _2099_ (.A(net72),
    .B_N(_0371_),
    .Y(\counter_lo_i.s_count [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2100_ (.Y(_0372_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(net5),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2101_ (.A(wdata_i[2]),
    .B(net67),
    .Y(_0373_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2102_ (.VSS(VSS),
    .VDD(VDD),
    .A1(net67),
    .A2(_0372_),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_nor2b_1 _2103_ (.A(net72),
    .B_N(_0374_),
    .Y(\counter_lo_i.s_count [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2104_ (.A(wdata_i[28]),
    .B(net64),
    .Y(_0375_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2105_ (.Y(_0376_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .B(_0270_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2106_ (.A(_0255_),
    .B(net19),
    .C(_0376_),
    .Y(_0377_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2107_ (.B(_0377_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .X(_0378_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2108_ (.A(net94),
    .B(_0378_),
    .Y(_0379_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2109_ (.A(net69),
    .B(_0375_),
    .C(_0379_),
    .Y(\counter_lo_i.s_count [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2110_ (.A(wdata_i[1]),
    .B(net67),
    .Y(_0380_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2111_ (.B(_1000_),
    .C(_0259_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .Y(_0381_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2112_ (.Y(_0382_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .B(_0381_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2113_ (.A(net95),
    .B(_0382_),
    .Y(_0383_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2114_ (.A(net72),
    .B(_0380_),
    .C(_0383_),
    .Y(\counter_lo_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2115_ (.A(wdata_i[0]),
    .B(net67),
    .Y(_0384_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2116_ (.Y(_0385_),
    .A(_1000_),
    .B(_0259_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2117_ (.A0(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_A ),
    .A1(\counter_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .S(_0385_),
    .X(_0386_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2118_ (.A(net95),
    .B(_0386_),
    .Y(_0387_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2119_ (.A(net72),
    .B(_0384_),
    .C(_0387_),
    .Y(\counter_lo_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2120_ (.A(wdata_i[27]),
    .B(net66),
    .Y(_0388_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2121_ (.VDD(VDD),
    .Y(_0389_),
    .A(_0270_),
    .VSS(VSS));
 sg13g2_nor3_1 _2122_ (.A(_0255_),
    .B(net19),
    .C(_0389_),
    .Y(_0390_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2123_ (.B(_0390_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .X(_0391_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2124_ (.A(net94),
    .B(_0391_),
    .Y(_0392_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2125_ (.A(net69),
    .B(_0388_),
    .C(_0392_),
    .Y(\counter_lo_i.s_count [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2126_ (.A(wdata_i[26]),
    .B(net65),
    .Y(_0393_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _2127_ (.A(_0255_),
    .B(net19),
    .C(_0269_),
    .Y(_0394_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _2128_ (.A(_0266_),
    .B_N(_0394_),
    .Y(_0395_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2129_ (.Y(_0396_),
    .A(_0265_),
    .B(_0395_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2130_ (.A(net93),
    .B(_0396_),
    .Y(_0397_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2131_ (.A(net70),
    .B(_0393_),
    .C(_0397_),
    .Y(\counter_lo_i.s_count [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2132_ (.A(wdata_i[25]),
    .B(net64),
    .Y(_0398_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2133_ (.Y(_0399_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .B(_0394_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2134_ (.Y(_0400_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .B(_0399_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2135_ (.A(net94),
    .B(_0400_),
    .Y(_0401_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2136_ (.A(net69),
    .B(_0398_),
    .C(_0401_),
    .Y(\counter_lo_i.s_count [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2137_ (.A(wdata_i[24]),
    .B(net65),
    .Y(_0402_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2138_ (.VDD(VDD),
    .Y(_0403_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .VSS(VSS));
 sg13g2_xnor2_1 _2139_ (.Y(_0404_),
    .A(_0403_),
    .B(_0394_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2140_ (.A(net93),
    .B(_0404_),
    .Y(_0405_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2141_ (.A(net70),
    .B(_0402_),
    .C(_0405_),
    .Y(\counter_lo_i.s_count [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2142_ (.A(wdata_i[23]),
    .B(net64),
    .Y(_0406_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _2143_ (.X(_0407_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(\counter_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .C(_0284_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2144_ (.B(_0407_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .X(_0408_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2145_ (.A(net94),
    .B(_0408_),
    .Y(_0409_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2146_ (.A(net69),
    .B(_0406_),
    .C(_0409_),
    .Y(\counter_lo_i.s_count [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2147_ (.A(wdata_i[22]),
    .B(net64),
    .Y(_0410_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2148_ (.Y(_0411_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .B(_0284_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2149_ (.Y(_0412_),
    .A(\counter_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(_0411_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2150_ (.A(net94),
    .B(_0412_),
    .Y(_0413_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2151_ (.A(net69),
    .B(_0410_),
    .C(_0413_),
    .Y(\counter_lo_i.s_count [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2152_ (.Y(_0414_),
    .A(\counter_lo_i.compare_value_i [20]),
    .B(\counter_lo_i.s_count [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2153_ (.Y(_0415_),
    .A(\counter_lo_i.compare_value_i [12]),
    .B(\counter_lo_i.s_count [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2154_ (.B(\counter_lo_i.s_count [8]),
    .A(\counter_lo_i.compare_value_i [8]),
    .X(_0416_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2155_ (.B(\counter_lo_i.s_count [6]),
    .A(\counter_lo_i.compare_value_i [6]),
    .X(_0417_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2156_ (.Y(_0418_),
    .A(\counter_lo_i.compare_value_i [2]),
    .B(\counter_lo_i.s_count [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2157_ (.Y(_0419_),
    .A(\counter_lo_i.compare_value_i [1]),
    .B(\counter_lo_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2158_ (.Y(_0420_),
    .A(\counter_lo_i.compare_value_i [4]),
    .B(\counter_lo_i.s_count [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2159_ (.Y(_0421_),
    .A(\counter_lo_i.compare_value_i [0]),
    .B(\counter_lo_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2160_ (.B(_0419_),
    .C(_0420_),
    .A(_0418_),
    .Y(_0422_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0421_));
 sg13g2_xnor2_1 _2161_ (.Y(_0423_),
    .A(\counter_lo_i.compare_value_i [7]),
    .B(\counter_lo_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2162_ (.Y(_0424_),
    .A(\counter_lo_i.compare_value_i [5]),
    .B(\counter_lo_i.s_count [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2163_ (.Y(_0425_),
    .A(_0423_),
    .B(_0424_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _2164_ (.A(_0416_),
    .B(_0417_),
    .C(_0422_),
    .Y(_0426_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0425_));
 sg13g2_xor2_1 _2165_ (.B(\counter_lo_i.s_count [16]),
    .A(\counter_lo_i.compare_value_i [16]),
    .X(_0427_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2166_ (.B(\counter_lo_i.s_count [15]),
    .A(\counter_lo_i.compare_value_i [15]),
    .X(_0428_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2167_ (.B(\counter_lo_i.s_count [18]),
    .A(\counter_lo_i.compare_value_i [18]),
    .X(_0429_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2168_ (.B(\counter_lo_i.s_count [17]),
    .A(\counter_lo_i.compare_value_i [17]),
    .X(_0430_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2169_ (.A(_0427_),
    .B(_0428_),
    .C(_0429_),
    .D(_0430_),
    .Y(_0431_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2170_ (.B(_0415_),
    .C(_0426_),
    .A(_0414_),
    .Y(_0432_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0431_));
 sg13g2_xnor2_1 _2171_ (.Y(_0433_),
    .A(\counter_lo_i.compare_value_i [26]),
    .B(\counter_lo_i.s_count [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2172_ (.B(\counter_lo_i.s_count [10]),
    .A(\counter_lo_i.compare_value_i [10]),
    .X(_0434_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2173_ (.B(\counter_lo_i.s_count [14]),
    .A(\counter_lo_i.compare_value_i [14]),
    .X(_0435_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2174_ (.B(\counter_lo_i.s_count [13]),
    .A(\counter_lo_i.compare_value_i [13]),
    .X(_0436_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2175_ (.B(\counter_lo_i.s_count [11]),
    .A(\counter_lo_i.compare_value_i [11]),
    .X(_0437_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _2176_ (.A(_0434_),
    .B(_0435_),
    .C(_0436_),
    .Y(_0438_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0437_));
 sg13g2_nand2_1 _2177_ (.Y(_0439_),
    .A(_0433_),
    .B(_0438_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2178_ (.Y(_0440_),
    .A(\counter_lo_i.compare_value_i [30]),
    .B(\counter_lo_i.s_count [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2179_ (.Y(_0441_),
    .A(\counter_lo_i.compare_value_i [25]),
    .B(\counter_lo_i.s_count [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2180_ (.Y(_0442_),
    .A(\counter_lo_i.compare_value_i [22]),
    .B(\counter_lo_i.s_count [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2181_ (.Y(_0443_),
    .A(\counter_lo_i.compare_value_i [23]),
    .B(\counter_lo_i.s_count [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2182_ (.B(_0441_),
    .C(_0442_),
    .A(_0440_),
    .Y(_0444_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0443_));
 sg13g2_xnor2_1 _2183_ (.Y(_0445_),
    .A(\counter_lo_i.compare_value_i [31]),
    .B(\counter_lo_i.s_count [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2184_ (.Y(_0446_),
    .A(\counter_lo_i.compare_value_i [24]),
    .B(\counter_lo_i.s_count [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2185_ (.B(\counter_lo_i.s_count [28]),
    .A(\counter_lo_i.compare_value_i [28]),
    .X(_0447_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2186_ (.B(\counter_lo_i.s_count [21]),
    .A(\counter_lo_i.compare_value_i [21]),
    .X(_0448_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2187_ (.A(_0447_),
    .B(_0448_),
    .Y(_0449_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2188_ (.A0(wdata_i[9]),
    .A1(_0343_),
    .S(net68),
    .X(_0450_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2189_ (.VDD(VDD),
    .Y(_0451_),
    .A(\counter_lo_i.compare_value_i [3]),
    .VSS(VSS));
 sg13g2_nand3_1 _2190_ (.B(_0366_),
    .C(_0370_),
    .A(_0451_),
    .Y(_0452_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21o_1 _2191_ (.A2(_0370_),
    .A1(_0366_),
    .B1(_0451_),
    .X(_0453_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2192_ (.B(_0450_),
    .C(_0452_),
    .A(\counter_lo_i.compare_value_i [9]),
    .Y(_0454_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0453_));
 sg13g2_inv_1 _2193_ (.VDD(VDD),
    .Y(_0455_),
    .A(\counter_lo_i.compare_value_i [9]),
    .VSS(VSS));
 sg13g2_nand4_1 _2194_ (.B(_0455_),
    .C(_0345_),
    .A(\counter_lo_i.compare_value_i [3]),
    .Y(_0456_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0371_));
 sg13g2_and2_1 _2195_ (.A(_0454_),
    .B(_0456_),
    .X(_0457_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2196_ (.A(_0450_),
    .B(_0371_),
    .Y(_0458_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2197_ (.A(\counter_lo_i.compare_value_i [3]),
    .B(\counter_lo_i.compare_value_i [9]),
    .Y(_0459_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2198_ (.B1(_0459_),
    .VDD(VDD),
    .Y(_0460_),
    .VSS(VSS),
    .A1(net73),
    .A2(_0458_));
 sg13g2_o21ai_1 _2199_ (.B1(_0460_),
    .VDD(VDD),
    .Y(_0461_),
    .VSS(VSS),
    .A1(net72),
    .A2(_0457_));
 sg13g2_xnor2_1 _2200_ (.Y(_0462_),
    .A(\counter_lo_i.compare_value_i [27]),
    .B(\counter_lo_i.s_count [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2201_ (.Y(_0463_),
    .A(\counter_lo_i.compare_value_i [29]),
    .B(\counter_lo_i.s_count [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2202_ (.Y(_0464_),
    .A(\counter_lo_i.compare_value_i [19]),
    .B(\counter_lo_i.s_count [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _2203_ (.A(_0461_),
    .B(_0462_),
    .C(_0463_),
    .D(_0464_),
    .X(_0465_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2204_ (.B(_0446_),
    .C(_0449_),
    .A(_0445_),
    .Y(_0466_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0465_));
 sg13g2_nor4_1 _2205_ (.A(_0432_),
    .B(_0439_),
    .C(_0444_),
    .D(_0466_),
    .Y(\counter_lo_i.target_reached_o_reg_D ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2206_ (.Y(_0467_),
    .A(_0941_),
    .B(_1140_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2207_ (.A0(wdata_i[3]),
    .A1(s_cfg_hi_reg[3]),
    .S(net90),
    .X(s_cfg_hi[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_2 _2208_ (.A(_1140_),
    .B(_0229_),
    .X(_0468_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net43),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2210_ (.A0(s_cfg_lo_reg[3]),
    .A1(wdata_i[3]),
    .S(net84),
    .X(s_cfg_lo[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_2 _2211_ (.X(irq_hi_o),
    .A(_0238_),
    .B(\counter_hi_i.target_reached_o ),
    .C(s_cfg_hi_reg[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2212_ (.VDD(VDD),
    .Y(_0470_),
    .A(s_cfg_lo_reg[2]),
    .VSS(VSS));
 sg13g2_nor2_2 _2213_ (.A(_0470_),
    .B(_0239_),
    .Y(irq_lo_o),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(net43),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2215_ (.A0(wdata_i[8]),
    .A1(\prescaler_hi_i.compare_value_i [0]),
    .S(net92),
    .X(_0064_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2216_ (.A0(wdata_i[9]),
    .A1(\prescaler_hi_i.compare_value_i [1]),
    .S(net91),
    .X(_0065_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2217_ (.A0(wdata_i[10]),
    .A1(\prescaler_hi_i.compare_value_i [2]),
    .S(net91),
    .X(_0066_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2218_ (.A0(wdata_i[11]),
    .A1(\prescaler_hi_i.compare_value_i [3]),
    .S(net91),
    .X(_0067_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2219_ (.A0(wdata_i[12]),
    .A1(\prescaler_hi_i.compare_value_i [4]),
    .S(net91),
    .X(_0068_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2220_ (.A0(wdata_i[13]),
    .A1(\prescaler_hi_i.compare_value_i [5]),
    .S(net91),
    .X(_0069_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2221_ (.A0(wdata_i[14]),
    .A1(\prescaler_hi_i.compare_value_i [6]),
    .S(net91),
    .X(_0070_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(net43),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2223_ (.A0(wdata_i[15]),
    .A1(\prescaler_hi_i.compare_value_i [7]),
    .S(net89),
    .X(_0071_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _2224_ (.B(_0953_),
    .C(_0959_),
    .Y(_0473_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\prescaler_hi_i.target_reached_o ));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(net43),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2226_ (.A(s_cfg_hi_reg[6]),
    .B(s_cfg_hi_reg[7]),
    .X(_0475_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _2227_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0476_),
    .B(\prescaler_hi_i.enable_count_i_$_AND__Y_B_$_MUX__Y_S_$_AND__Y_B ),
    .A(s_cfg_hi_reg[7]));
 sg13g2_a221oi_1 _2228_ (.VSS(VSS),
    .VDD(VDD),
    .B2(\prescaler_hi_i.target_reached_o_$_MUX__A_S_$_AND__Y_A ),
    .C1(_0934_),
    .B1(_0476_),
    .A1(_0978_),
    .Y(_0477_),
    .A2(_0475_));
 sg13g2_and3_1 _2229_ (.X(_0478_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _2230_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .C(_0477_),
    .D(_0478_),
    .X(_0479_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2231_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .B(_0479_),
    .X(_0480_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2232_ (.Y(_0481_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(_0480_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2233_ (.B(_0481_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .X(_0482_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2234_ (.A(net78),
    .B(_0482_),
    .Y(\prescaler_hi_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2235_ (.Y(_0483_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(_0480_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2236_ (.A(net78),
    .B(_0483_),
    .Y(\prescaler_hi_i.s_count [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2237_ (.Y(_0484_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .B(_0479_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2238_ (.A(net77),
    .B(_0484_),
    .Y(\prescaler_hi_i.s_count [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2239_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .B(_0477_),
    .X(_0485_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2240_ (.Y(_0486_),
    .A(_0485_),
    .B(_0478_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2241_ (.B(_0486_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .X(_0487_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2242_ (.A(net77),
    .B(_0487_),
    .Y(\prescaler_hi_i.s_count [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2243_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .C(_0485_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .Y(_0488_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2244_ (.B(_0488_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .X(_0489_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2245_ (.A(net77),
    .B(_0489_),
    .Y(\prescaler_hi_i.s_count [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2246_ (.Y(_0490_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .B(_0485_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2247_ (.B(_0490_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .X(_0491_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2248_ (.A(net77),
    .B(_0491_),
    .Y(\prescaler_hi_i.s_count [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2249_ (.Y(_0492_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .B(_0485_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2250_ (.A(net77),
    .B(_0492_),
    .Y(\prescaler_hi_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _2251_ (.Y(_0493_),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .A_N(_0477_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2252_ (.Y(_0494_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [0]),
    .B(_0477_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2253_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_0493_),
    .A2(_0494_),
    .Y(\prescaler_hi_i.s_count [0]),
    .B1(net77));
 sg13g2_buf_2 fanout38 (.A(_0742_),
    .X(net38),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2255_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .Y(_0496_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]));
 sg13g2_inv_1 _2256_ (.VDD(VDD),
    .Y(_0497_),
    .A(_0496_),
    .VSS(VSS));
 sg13g2_inv_1 _2257_ (.VDD(VDD),
    .Y(_0498_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .VSS(VSS));
 sg13g2_inv_2 _2258_ (.Y(_0499_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2259_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .X(_0500_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2260_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .C(_0479_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .Y(_0501_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0500_));
 sg13g2_nand3_1 _2261_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .Y(_0502_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2262_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .Y(_0503_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [14]));
 sg13g2_nor2_1 _2263_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2264_ (.Y(_0505_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .B(_0504_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_2 _2265_ (.A(_0498_),
    .B(_0499_),
    .C(_0501_),
    .Y(_0506_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0505_));
 sg13g2_and4_2 _2266_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .D(_0506_),
    .X(_0507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout37 (.A(net38),
    .X(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _2268_ (.X(_0509_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .B(_0497_),
    .C(_0507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _2269_ (.X(_0510_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .C(_0509_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2270_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .C(_0510_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .Y(_0511_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2271_ (.B(_0511_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .X(_0512_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2272_ (.A(net79),
    .B(_0512_),
    .Y(\prescaler_hi_i.s_count [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2273_ (.Y(_0513_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .B(_0510_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2274_ (.B(_0513_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .X(_0514_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2275_ (.A(net79),
    .B(_0514_),
    .Y(\prescaler_hi_i.s_count [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2276_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .B(_0506_),
    .X(_0515_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2277_ (.Y(_0516_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(_0515_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2278_ (.B(_0516_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .X(_0517_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2279_ (.A(net81),
    .B(_0517_),
    .Y(\prescaler_hi_i.s_count [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2280_ (.Y(_0518_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(_0515_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2281_ (.A(net80),
    .B(_0518_),
    .Y(\prescaler_hi_i.s_count [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2282_ (.Y(_0519_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .B(_0506_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2283_ (.A(net80),
    .B(_0519_),
    .Y(\prescaler_hi_i.s_count [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_2 _2284_ (.A(_0498_),
    .B(_0499_),
    .C(_0501_),
    .Y(_0520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2285_ (.Y(_0521_),
    .A(_0504_),
    .B(_0520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2286_ (.B(_0521_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .X(_0522_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2287_ (.A(net80),
    .B(_0522_),
    .Y(\prescaler_hi_i.s_count [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2288_ (.VDD(VDD),
    .Y(_0523_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .VSS(VSS));
 sg13g2_inv_1 _2289_ (.VDD(VDD),
    .Y(_0524_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .VSS(VSS));
 sg13g2_nand2b_2 _2290_ (.Y(_0525_),
    .B(_0520_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(_0502_));
 sg13g2_nor3_1 _2291_ (.A(_0523_),
    .B(_0524_),
    .C(_0525_),
    .Y(_0526_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2292_ (.Y(_0527_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .B(_0526_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2293_ (.B(_0527_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .X(_0528_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2294_ (.A(net80),
    .B(_0528_),
    .Y(\prescaler_hi_i.s_count [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2295_ (.Y(_0529_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .B(_0526_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2296_ (.A(net80),
    .B(_0529_),
    .Y(\prescaler_hi_i.s_count [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2297_ (.A(_0524_),
    .B(_0525_),
    .Y(_0530_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2298_ (.Y(_0531_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .B(_0530_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2299_ (.A(net80),
    .B(_0531_),
    .Y(\prescaler_hi_i.s_count [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout36 (.A(net38),
    .X(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2301_ (.Y(_0533_),
    .A(_0524_),
    .B(_0525_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2302_ (.A(net81),
    .B(_0533_),
    .Y(\prescaler_hi_i.s_count [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2303_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .C(_0520_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .Y(_0534_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2304_ (.B(_0534_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .X(_0535_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2305_ (.A(net78),
    .B(_0535_),
    .Y(\prescaler_hi_i.s_count [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2306_ (.Y(_0536_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .B(_0520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2307_ (.B(_0536_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .X(_0537_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2308_ (.A(net80),
    .B(_0537_),
    .Y(\prescaler_hi_i.s_count [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2309_ (.Y(_0538_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .B(_0510_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2310_ (.A(net79),
    .B(_0538_),
    .Y(\prescaler_hi_i.s_count [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2311_ (.Y(_0539_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .B(_0520_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2312_ (.A(net78),
    .B(_0539_),
    .Y(\prescaler_hi_i.s_count [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2313_ (.A(_0499_),
    .B(_0501_),
    .Y(_0540_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2314_ (.Y(_0541_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(_0540_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2315_ (.A(net80),
    .B(_0541_),
    .Y(\prescaler_hi_i.s_count [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2316_ (.Y(_0542_),
    .A(_0499_),
    .B(_0501_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2317_ (.A(net77),
    .B(_0542_),
    .Y(\prescaler_hi_i.s_count [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2318_ (.Y(_0543_),
    .A(_0480_),
    .B(_0500_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2319_ (.Y(_0544_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(_0543_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _2320_ (.A(net77),
    .B_N(_0544_),
    .Y(\prescaler_hi_i.s_count [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2321_ (.Y(_0545_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .B(_0509_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2322_ (.B(_0545_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .X(_0546_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2323_ (.A(net79),
    .B(_0546_),
    .Y(\prescaler_hi_i.s_count [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2324_ (.Y(_0547_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .B(_0509_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2325_ (.A(net81),
    .B(_0547_),
    .Y(\prescaler_hi_i.s_count [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2326_ (.Y(_0548_),
    .A(_0497_),
    .B(_0507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2327_ (.B(_0548_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .X(_0549_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2328_ (.A(net81),
    .B(_0549_),
    .Y(\prescaler_hi_i.s_count [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2329_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .Y(_0550_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0507_));
 sg13g2_xor2_1 _2330_ (.B(_0550_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .X(_0551_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2331_ (.A(net79),
    .B(_0551_),
    .Y(\prescaler_hi_i.s_count [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2332_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .C(_0507_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .Y(_0552_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2333_ (.B(_0552_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .X(_0553_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2334_ (.A(net79),
    .B(_0553_),
    .Y(\prescaler_hi_i.s_count [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2335_ (.Y(_0554_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(_0507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2336_ (.B(_0554_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .X(_0555_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2337_ (.A(net79),
    .B(_0555_),
    .Y(\prescaler_hi_i.s_count [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2338_ (.Y(_0556_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(_0507_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2339_ (.A(net79),
    .B(_0556_),
    .Y(\prescaler_hi_i.s_count [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_1 _2340_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .X(_0557_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 _2341_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .C(_0509_),
    .D(_0557_),
    .X(_0558_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2342_ (.B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .Y(_0559_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0510_));
 sg13g2_nand3_1 _2343_ (.B(_0497_),
    .C(_0507_),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .Y(_0560_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2344_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .D(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .Y(_0561_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2345_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .D(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .Y(_0562_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _2346_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0563_),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [26]));
 sg13g2_nor4_1 _2347_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .D(_0563_),
    .Y(_0564_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2348_ (.B(_0561_),
    .C(_0562_),
    .A(_0525_),
    .Y(_0565_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0564_));
 sg13g2_nand2_1 _2349_ (.Y(_0566_),
    .A(_0498_),
    .B(_0499_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2350_ (.A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .C(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .D(_0566_),
    .Y(_0567_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _2351_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0568_),
    .B(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .A(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [12]));
 sg13g2_o21ai_1 _2352_ (.B1(_0502_),
    .VDD(VDD),
    .Y(_0569_),
    .VSS(VSS),
    .A1(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .A2(_0568_));
 sg13g2_a22oi_1 _2353_ (.Y(_0570_),
    .B1(_0569_),
    .B2(_0520_),
    .A2(_0567_),
    .A1(_0543_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a221oi_1 _2354_ (.VSS(VSS),
    .VDD(VDD),
    .B2(_0565_),
    .C1(_0570_),
    .B1(_0560_),
    .A1(_0558_),
    .Y(_0571_),
    .A2(_0559_));
 sg13g2_nor2_1 _2355_ (.A(net78),
    .B(_0571_),
    .Y(_0572_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2356_ (.Y(_0573_),
    .A(\prescaler_hi_i.compare_value_i [6]),
    .B(\prescaler_hi_i.s_count [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2357_ (.Y(_0574_),
    .A(\prescaler_hi_i.compare_value_i [7]),
    .B(\prescaler_hi_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2358_ (.B(\prescaler_hi_i.s_count [4]),
    .A(\prescaler_hi_i.compare_value_i [4]),
    .X(_0575_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2359_ (.B(\prescaler_hi_i.s_count [3]),
    .A(\prescaler_hi_i.compare_value_i [3]),
    .X(_0576_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2360_ (.B(\prescaler_hi_i.s_count [5]),
    .A(\prescaler_hi_i.compare_value_i [5]),
    .X(_0577_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2361_ (.Y(_0578_),
    .A(\prescaler_hi_i.compare_value_i [2]),
    .B(\prescaler_hi_i.s_count [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2362_ (.Y(_0579_),
    .A(\prescaler_hi_i.compare_value_i [0]),
    .B(\prescaler_hi_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2363_ (.Y(_0580_),
    .A(\prescaler_hi_i.compare_value_i [1]),
    .B(\prescaler_hi_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2364_ (.B(_0579_),
    .C(_0580_),
    .A(_0578_),
    .Y(_0581_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2365_ (.A(_0575_),
    .B(_0576_),
    .C(_0577_),
    .D(_0581_),
    .Y(_0582_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2366_ (.B(_0574_),
    .C(_0582_),
    .A(_0573_),
    .Y(_0583_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2367_ (.A(\prescaler_hi_i.s_count [11]),
    .B(_0572_),
    .C(_0583_),
    .Y(\prescaler_hi_i.target_reached_o_reg_D ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout35 (.A(net38),
    .X(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2369_ (.A0(\prescaler_lo_i.compare_value_i [0]),
    .A1(wdata_i[8]),
    .S(net86),
    .X(_0072_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2370_ (.A0(\prescaler_lo_i.compare_value_i [1]),
    .A1(wdata_i[9]),
    .S(net86),
    .X(_0073_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout34 (.A(net38),
    .X(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2372_ (.VDD(VDD),
    .Y(_0586_),
    .A(\prescaler_lo_i.compare_value_i [2]),
    .VSS(VSS));
 sg13g2_buf_2 fanout33 (.A(_0743_),
    .X(net33),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2374_ (.Y(_0588_),
    .A(wdata_i[10]),
    .B(net87),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2375_ (.B1(_0588_),
    .VDD(VDD),
    .Y(_0074_),
    .VSS(VSS),
    .A1(_0586_),
    .A2(net87));
 sg13g2_mux2_1 _2376_ (.A0(\prescaler_lo_i.compare_value_i [3]),
    .A1(wdata_i[11]),
    .S(net86),
    .X(_0075_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2377_ (.A0(\prescaler_lo_i.compare_value_i [4]),
    .A1(wdata_i[12]),
    .S(net86),
    .X(_0076_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2378_ (.A0(\prescaler_lo_i.compare_value_i [5]),
    .A1(wdata_i[13]),
    .S(net86),
    .X(_0077_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2379_ (.A0(\prescaler_lo_i.compare_value_i [6]),
    .A1(wdata_i[14]),
    .S(net86),
    .X(_0078_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2380_ (.A0(\prescaler_lo_i.compare_value_i [7]),
    .A1(wdata_i[15]),
    .S(net83),
    .X(_0079_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2381_ (.Y(_0589_),
    .A(_0998_),
    .B(_0241_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2382_ (.VDD(VDD),
    .Y(_0590_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .VSS(VSS));
 sg13g2_buf_2 fanout32 (.A(net33),
    .X(net32),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout31 (.A(net32),
    .X(net31),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2385_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .X(_0593_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2386_ (.VDD(VDD),
    .Y(_0594_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .VSS(VSS));
 sg13g2_inv_1 _2387_ (.VDD(VDD),
    .Y(_0595_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .VSS(VSS));
 sg13g2_a21oi_1 _2388_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ),
    .A2(\counter_lo_i.enable_count_i_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_B ),
    .Y(_0596_),
    .B1(s_cfg_lo_reg[7]));
 sg13g2_a21oi_1 _2389_ (.VSS(VSS),
    .VDD(VDD),
    .A1(s_cfg_lo_reg[6]),
    .A2(_0978_),
    .Y(_0597_),
    .B1(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ));
 sg13g2_o21ai_1 _2390_ (.B1(s_cfg_lo_reg[0]),
    .VDD(VDD),
    .Y(_0598_),
    .VSS(VSS),
    .A1(_0596_),
    .A2(_0597_));
 sg13g2_nor3_2 _2391_ (.A(_0594_),
    .B(_0595_),
    .C(_0598_),
    .Y(_0599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _2392_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .C(_0593_),
    .D(_0599_),
    .X(_0600_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_2 _2393_ (.Y(_0601_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(_0600_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2394_ (.Y(_0602_),
    .A(_0590_),
    .B(_0601_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2395_ (.A(net60),
    .B(_0602_),
    .Y(\prescaler_lo_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout30 (.A(net33),
    .X(net30),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2397_ (.Y(_0604_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .B(_0600_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2398_ (.A(net62),
    .B(_0604_),
    .Y(\prescaler_lo_i.s_count [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2399_ (.B(_0593_),
    .C(_0599_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .Y(_0605_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2400_ (.B(_0605_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .X(_0606_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2401_ (.A(net62),
    .B(_0606_),
    .Y(\prescaler_lo_i.s_count [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2402_ (.Y(_0607_),
    .A(_0593_),
    .B(_0599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2403_ (.B(_0607_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .X(_0608_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2404_ (.A(net62),
    .B(_0608_),
    .Y(\prescaler_lo_i.s_count [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout29 (.A(net33),
    .X(net29),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2406_ (.Y(_0610_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(_0599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2407_ (.B(_0610_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .X(_0611_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2408_ (.A(net62),
    .B(_0611_),
    .Y(\prescaler_lo_i.s_count [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2409_ (.Y(_0612_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(_0599_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2410_ (.A(net62),
    .B(_0612_),
    .Y(\prescaler_lo_i.s_count [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2411_ (.A(_0595_),
    .B(_0598_),
    .Y(_0613_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2412_ (.Y(_0614_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .B(_0613_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2413_ (.A(net62),
    .B(_0614_),
    .Y(\prescaler_lo_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2414_ (.A(_0998_),
    .B(_0241_),
    .X(_0615_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2415_ (.A0(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [0]),
    .A1(\prescaler_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .S(_0598_),
    .X(_0616_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2416_ (.A(_0615_),
    .B(_0616_),
    .X(\prescaler_lo_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2417_ (.VDD(VDD),
    .Y(_0617_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [31]),
    .VSS(VSS));
 sg13g2_inv_1 _2418_ (.VDD(VDD),
    .Y(_0618_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .VSS(VSS));
 sg13g2_inv_1 _2419_ (.VDD(VDD),
    .Y(_0619_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .VSS(VSS));
 sg13g2_nand2_1 _2420_ (.Y(_0620_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2421_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .X(_0621_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _2422_ (.X(_0622_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _2423_ (.X(_0623_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _2424_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .C(_0622_),
    .D(_0623_),
    .X(_0624_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2425_ (.B(_0621_),
    .C(_0624_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .Y(_0625_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2426_ (.A(_0619_),
    .B(_0620_),
    .C(_0625_),
    .Y(_0626_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _2427_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .D(_0626_),
    .X(_0627_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2428_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .C(_0600_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .Y(_0628_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0627_));
 sg13g2_nand3_1 _2429_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .Y(_0629_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2430_ (.A(_0618_),
    .B(_0628_),
    .C(_0629_),
    .Y(_0630_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2431_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .B(_0630_),
    .X(_0631_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2432_ (.Y(_0632_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .B(_0631_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2433_ (.Y(_0633_),
    .A(_0617_),
    .B(_0632_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2434_ (.A(net61),
    .B(_0633_),
    .Y(\prescaler_lo_i.s_count [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2435_ (.Y(_0634_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .B(_0631_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2436_ (.A(net61),
    .B(_0634_),
    .Y(\prescaler_lo_i.s_count [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_2 _2437_ (.A(_0601_),
    .B_N(_0626_),
    .Y(_0635_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2438_ (.Y(_0636_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .B(_0635_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2439_ (.A(net61),
    .B(_0636_),
    .Y(\prescaler_lo_i.s_count [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _2440_ (.A(_0601_),
    .B(_0625_),
    .Y(_0637_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2441_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .C(_0637_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .Y(_0638_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2442_ (.B(_0638_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .X(_0639_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2443_ (.A(net60),
    .B(_0639_),
    .Y(\prescaler_lo_i.s_count [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2444_ (.Y(_0640_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .B(_0637_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2445_ (.B(_0640_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .X(_0641_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2446_ (.A(net59),
    .B(_0641_),
    .Y(\prescaler_lo_i.s_count [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2447_ (.Y(_0642_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .B(_0637_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2448_ (.A(net59),
    .B(_0642_),
    .Y(\prescaler_lo_i.s_count [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _2449_ (.A(_0590_),
    .B(_0601_),
    .Y(_0643_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2450_ (.B(_0624_),
    .C(_0643_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .Y(_0644_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2451_ (.B(_0644_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .X(_0645_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2452_ (.A(net60),
    .B(_0645_),
    .Y(\prescaler_lo_i.s_count [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2453_ (.Y(_0646_),
    .A(_0624_),
    .B(_0643_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2454_ (.B(_0646_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .X(_0647_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2455_ (.A(net59),
    .B(_0647_),
    .Y(\prescaler_lo_i.s_count [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout28 (.X(net28),
    .A(_1005_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_2 _2457_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .C(_0622_),
    .D(_0643_),
    .X(_0649_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2458_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .C(_0649_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .Y(_0650_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2459_ (.B(_0650_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .X(_0651_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2460_ (.A(net59),
    .B(_0651_),
    .Y(\prescaler_lo_i.s_count [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2461_ (.Y(_0652_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .B(_0649_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2462_ (.B(_0652_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .X(_0653_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2463_ (.A(net59),
    .B(_0653_),
    .Y(\prescaler_lo_i.s_count [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2464_ (.Y(_0654_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .B(_0649_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2465_ (.A(net59),
    .B(_0654_),
    .Y(\prescaler_lo_i.s_count [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2466_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .Y(_0655_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_2 _2467_ (.A(_0601_),
    .B(_0655_),
    .Y(_0656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _2468_ (.X(_0657_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .C(_0656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2469_ (.Y(_0658_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .B(_0657_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2470_ (.A(net59),
    .B(_0658_),
    .Y(\prescaler_lo_i.s_count [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2471_ (.Y(_0659_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .B(_0630_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2472_ (.A(net63),
    .B(_0659_),
    .Y(\prescaler_lo_i.s_count [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2473_ (.Y(_0660_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(_0656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2474_ (.B(_0660_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .X(_0661_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2475_ (.A(net59),
    .B(_0661_),
    .Y(\prescaler_lo_i.s_count [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2476_ (.Y(_0662_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(_0656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2477_ (.A(net60),
    .B(_0662_),
    .Y(\prescaler_lo_i.s_count [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2478_ (.Y(_0663_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(_0643_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2479_ (.B(_0663_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .X(_0664_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2480_ (.A(net60),
    .B(_0664_),
    .Y(\prescaler_lo_i.s_count [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2481_ (.Y(_0665_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(_0643_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2482_ (.A(net60),
    .B(_0665_),
    .Y(\prescaler_lo_i.s_count [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2483_ (.A(_0618_),
    .B(_0628_),
    .Y(_0666_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2484_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .C(_0666_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .Y(_0667_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2485_ (.B(_0667_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .X(_0668_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2486_ (.A(net63),
    .B(_0668_),
    .Y(\prescaler_lo_i.s_count [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2487_ (.Y(_0669_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .B(_0666_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2488_ (.B(_0669_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .X(_0670_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2489_ (.A(net61),
    .B(_0670_),
    .Y(\prescaler_lo_i.s_count [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2490_ (.Y(_0671_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .B(_0666_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2491_ (.A(net61),
    .B(_0671_),
    .Y(\prescaler_lo_i.s_count [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2492_ (.Y(_0672_),
    .A(_0618_),
    .B(_0628_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2493_ (.A(net61),
    .B(_0672_),
    .Y(\prescaler_lo_i.s_count [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _2494_ (.A(_0601_),
    .B_N(_0627_),
    .Y(_0673_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2495_ (.Y(_0674_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .B(_0673_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2496_ (.A(net62),
    .B(_0674_),
    .Y(\prescaler_lo_i.s_count [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2497_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .C(_0635_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .Y(_0675_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2498_ (.B(_0675_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .X(_0676_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2499_ (.A(net61),
    .B(_0676_),
    .Y(\prescaler_lo_i.s_count [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2500_ (.Y(_0677_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .B(_0635_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2501_ (.B(_0677_),
    .A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .X(_0678_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2502_ (.A(net61),
    .B(_0678_),
    .Y(\prescaler_lo_i.s_count [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 _2503_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .D(_0637_),
    .X(_0679_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2504_ (.B1(_0679_),
    .VDD(VDD),
    .Y(_0680_),
    .VSS(VSS),
    .A1(_0620_),
    .A2(_0640_));
 sg13g2_nor3_1 _2505_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [31]),
    .Y(_0681_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2506_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .D(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .Y(_0682_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2507_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .D(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .Y(_0683_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2508_ (.B(_0682_),
    .C(_0683_),
    .A(_0681_),
    .Y(_0684_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or2_1 _2509_ (.VSS(VSS),
    .VDD(VDD),
    .X(_0685_),
    .B(_0684_),
    .A(_0635_));
 sg13g2_o21ai_1 _2510_ (.B1(_0685_),
    .VDD(VDD),
    .Y(_0686_),
    .VSS(VSS),
    .A1(_0617_),
    .A2(_0632_));
 sg13g2_or4_1 _2511_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .D(_0656_),
    .X(_0687_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2512_ (.Y(_0688_),
    .A(_0622_),
    .B(_0656_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or4_1 _2513_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .D(_0649_),
    .X(_0689_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2514_ (.Y(_0690_),
    .A(_0623_),
    .B(_0649_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2515_ (.Y(_0691_),
    .B1(_0689_),
    .B2(_0690_),
    .A2(_0688_),
    .A1(_0687_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2516_ (.B(_0686_),
    .C(_0691_),
    .A(_0680_),
    .Y(_0692_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2517_ (.Y(_0693_),
    .A(\prescaler_lo_i.compare_value_i [6]),
    .B(\prescaler_lo_i.s_count [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2518_ (.Y(_0694_),
    .A(\prescaler_lo_i.compare_value_i [7]),
    .B(\prescaler_lo_i.s_count [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2519_ (.Y(_0695_),
    .A(\prescaler_lo_i.compare_value_i [2]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and2_1 _2520_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .B(_0695_),
    .X(_0696_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _2521_ (.Y(_0697_),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .A_N(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3b_1 _2522_ (.B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .C(\prescaler_lo_i.compare_value_i [2]),
    .Y(_0698_),
    .VDD(VDD),
    .VSS(VSS),
    .A_N(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]));
 sg13g2_o21ai_1 _2523_ (.B1(_0698_),
    .VDD(VDD),
    .Y(_0699_),
    .VSS(VSS),
    .A1(\prescaler_lo_i.compare_value_i [2]),
    .A2(_0697_));
 sg13g2_mux2_1 _2524_ (.A0(_0696_),
    .A1(_0699_),
    .S(_0599_),
    .X(_0700_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2525_ (.A(_0586_),
    .B(\prescaler_lo_i.compare_value_i [3]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .D(_0612_),
    .Y(_0701_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2526_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\prescaler_lo_i.compare_value_i [3]),
    .A2(_0700_),
    .Y(_0702_),
    .B1(_0701_));
 sg13g2_nor3_1 _2527_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .C(_0599_),
    .Y(_0703_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2528_ (.Y(_0704_),
    .A(_0615_),
    .B(_0607_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2529_ (.A(\prescaler_lo_i.compare_value_i [2]),
    .B(\prescaler_lo_i.compare_value_i [3]),
    .Y(_0705_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2530_ (.B1(_0705_),
    .VDD(VDD),
    .Y(_0706_),
    .VSS(VSS),
    .A1(_0703_),
    .A2(_0704_));
 sg13g2_o21ai_1 _2531_ (.B1(_0706_),
    .VDD(VDD),
    .Y(_0707_),
    .VSS(VSS),
    .A1(net62),
    .A2(_0702_));
 sg13g2_xnor2_1 _2532_ (.Y(_0708_),
    .A(\prescaler_lo_i.compare_value_i [4]),
    .B(\prescaler_lo_i.s_count [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2533_ (.Y(_0709_),
    .A(\prescaler_lo_i.compare_value_i [0]),
    .B(\prescaler_lo_i.s_count [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xnor2_1 _2534_ (.Y(_0710_),
    .A(\prescaler_lo_i.compare_value_i [1]),
    .B(\prescaler_lo_i.s_count [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and4_1 _2535_ (.A(_0707_),
    .B(_0708_),
    .C(_0709_),
    .D(_0710_),
    .X(_0711_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2536_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .C(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .D(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .Y(_0712_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2537_ (.B1(_0712_),
    .VDD(VDD),
    .Y(_0713_),
    .VSS(VSS),
    .A1(_0590_),
    .A2(_0601_));
 sg13g2_nor3_1 _2538_ (.A(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .B(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .C(_0624_),
    .Y(_0714_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2539_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_0621_),
    .A2(_0624_),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nor3_1 _2540_ (.A(_0601_),
    .B(_0655_),
    .C(_0715_),
    .Y(_0716_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2541_ (.A(net60),
    .B(_0716_),
    .Y(_0717_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_xor2_1 _2542_ (.B(\prescaler_lo_i.s_count [5]),
    .A(\prescaler_lo_i.compare_value_i [5]),
    .X(_0718_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2543_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_0713_),
    .A2(_0717_),
    .Y(_0719_),
    .B1(_0718_));
 sg13g2_nand4_1 _2544_ (.B(_0694_),
    .C(_0711_),
    .A(_0693_),
    .Y(_0720_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0719_));
 sg13g2_a21oi_1 _2545_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_0615_),
    .A2(_0692_),
    .Y(\prescaler_lo_i.target_reached_o_reg_D ),
    .B1(_0720_));
 sg13g2_buf_2 fanout27 (.A(net28),
    .X(net27),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2547_ (.VSS(VSS),
    .VDD(VDD),
    .A1(s_addr[4]),
    .A2(\s_addr_$_NOT__A_1_Y ),
    .Y(_0722_),
    .B1(s_addr[3]));
 sg13g2_nor2_1 _2548_ (.A(s_addr[4]),
    .B(\s_addr_$_NOT__A_Y ),
    .Y(_0723_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_or3_2 _2549_ (.A(s_addr[5]),
    .B(s_addr[0]),
    .C(s_addr[1]),
    .X(_0724_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout26 (.A(net27),
    .X(net26),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2551_ (.Y(_0726_),
    .A(s_addr[2]),
    .B(\s_addr_$_NOT__A_2_Y ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _2552_ (.B(s_wen),
    .C(_0726_),
    .A(r_valid_o),
    .Y(_0727_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2553_ (.A(_0724_),
    .B(_0727_),
    .Y(_0728_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2554_ (.B1(_0728_),
    .VDD(VDD),
    .Y(_0729_),
    .VSS(VSS),
    .A1(_0722_),
    .A2(_0723_));
 sg13g2_buf_2 fanout25 (.A(_0729_),
    .X(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2556_ (.A(s_addr[3]),
    .B(s_addr[4]),
    .C(\s_addr_$_NOT__A_2_Y ),
    .D(_0724_),
    .Y(_0731_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout24 (.X(net24),
    .A(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2558_ (.Y(_0733_),
    .A(s_cfg_hi_reg[31]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2559_ (.A(s_addr[3]),
    .B(s_addr[4]),
    .C(s_addr[2]),
    .D(_0724_),
    .Y(_0734_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(net24),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2561_ (.Y(_0736_),
    .A(s_cfg_lo_reg[31]),
    .B(net51),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2562_ (.A(s_addr[4]),
    .B(\s_addr_$_NOT__A_Y ),
    .C(\s_addr_$_NOT__A_2_Y ),
    .D(_0724_),
    .Y(_0737_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout22 (.X(net22),
    .A(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2564_ (.A(s_addr[4]),
    .B(s_addr[2]),
    .C(\s_addr_$_NOT__A_Y ),
    .D(_0724_),
    .Y(_0739_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout21 (.X(net21),
    .A(net25),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2566_ (.Y(_0741_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [31]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2567_ (.A(s_addr[3]),
    .B(s_addr[2]),
    .C(\s_addr_$_NOT__A_1_Y ),
    .D(_0724_),
    .Y(_0742_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _2568_ (.A(s_addr[3]),
    .B(\s_addr_$_NOT__A_2_Y ),
    .C(\s_addr_$_NOT__A_1_Y ),
    .D(_0724_),
    .Y(_0743_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout20 (.A(_0263_),
    .X(net20),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2570_ (.Y(_0745_),
    .B1(net31),
    .B2(\counter_hi_i.compare_value_i [31]),
    .A2(net37),
    .A1(\counter_lo_i.compare_value_i [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2571_ (.B(_0736_),
    .C(_0741_),
    .A(_0733_),
    .Y(_0746_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0745_));
 sg13g2_nor2b_2 _2572_ (.A(net23),
    .B_N(_0746_),
    .Y(r_rdata_o[31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2573_ (.Y(_0747_),
    .A(s_cfg_hi_reg[30]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout19 (.X(net19),
    .A(net20),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2575_ (.Y(_0749_),
    .A(\counter_lo_i.compare_value_i [30]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2576_ (.Y(_0750_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2577_ (.Y(_0751_),
    .B1(net49),
    .B2(s_cfg_lo_reg[30]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2578_ (.B(_0749_),
    .C(_0750_),
    .A(_0747_),
    .Y(_0752_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0751_));
 sg13g2_nor2b_2 _2579_ (.A(net22),
    .B_N(_0752_),
    .Y(r_rdata_o[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2580_ (.Y(_0753_),
    .A(s_cfg_hi_reg[21]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2581_ (.Y(_0754_),
    .A(\counter_lo_i.compare_value_i [21]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2582_ (.Y(_0755_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2583_ (.Y(_0756_),
    .B1(net49),
    .B2(s_cfg_lo_reg[21]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2584_ (.B(_0754_),
    .C(_0755_),
    .A(_0753_),
    .Y(_0757_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0756_));
 sg13g2_nor2b_2 _2585_ (.A(net21),
    .B_N(_0757_),
    .Y(r_rdata_o[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2586_ (.Y(_0758_),
    .A(s_cfg_hi_reg[20]),
    .B(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2587_ (.Y(_0759_),
    .A(\counter_lo_i.compare_value_i [20]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2588_ (.Y(_0760_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2589_ (.Y(_0761_),
    .B1(net50),
    .B2(s_cfg_lo_reg[20]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2590_ (.B(_0759_),
    .C(_0760_),
    .A(_0758_),
    .Y(_0762_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0761_));
 sg13g2_nor2b_2 _2591_ (.A(net22),
    .B_N(_0762_),
    .Y(r_rdata_o[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2592_ (.Y(_0763_),
    .A(s_cfg_hi_reg[19]),
    .B(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2593_ (.Y(_0764_),
    .A(\counter_lo_i.compare_value_i [19]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2594_ (.Y(_0765_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2595_ (.Y(_0766_),
    .B1(net50),
    .B2(s_cfg_lo_reg[19]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2596_ (.B(_0764_),
    .C(_0765_),
    .A(_0763_),
    .Y(_0767_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0766_));
 sg13g2_nor2b_2 _2597_ (.A(net21),
    .B_N(_0767_),
    .Y(r_rdata_o[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2598_ (.Y(_0768_),
    .A(s_cfg_hi_reg[18]),
    .B(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2599_ (.Y(_0769_),
    .A(\counter_lo_i.compare_value_i [18]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2600_ (.Y(_0770_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2601_ (.Y(_0771_),
    .B1(net50),
    .B2(s_cfg_lo_reg[18]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2602_ (.B(_0769_),
    .C(_0770_),
    .A(_0768_),
    .Y(_0772_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0771_));
 sg13g2_nor2b_2 _2603_ (.A(net21),
    .B_N(_0772_),
    .Y(r_rdata_o[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2604_ (.Y(_0773_),
    .A(s_cfg_hi_reg[17]),
    .B(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2605_ (.Y(_0774_),
    .A(\counter_lo_i.compare_value_i [17]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2606_ (.Y(_0775_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2607_ (.Y(_0776_),
    .B1(net50),
    .B2(s_cfg_lo_reg[17]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2608_ (.B(_0774_),
    .C(_0775_),
    .A(_0773_),
    .Y(_0777_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0776_));
 sg13g2_nor2b_2 _2609_ (.A(net22),
    .B_N(_0777_),
    .Y(r_rdata_o[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2610_ (.Y(_0778_),
    .A(s_cfg_hi_reg[16]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2611_ (.Y(_0779_),
    .A(\counter_lo_i.compare_value_i [16]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2612_ (.Y(_0780_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2613_ (.Y(_0781_),
    .B1(net51),
    .B2(s_cfg_lo_reg[16]),
    .A2(net31),
    .A1(\counter_hi_i.compare_value_i [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2614_ (.B(_0779_),
    .C(_0780_),
    .A(_0778_),
    .Y(_0782_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0781_));
 sg13g2_nor2b_2 _2615_ (.A(net23),
    .B_N(_0782_),
    .Y(r_rdata_o[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2616_ (.Y(_0783_),
    .A(\prescaler_hi_i.compare_value_i [7]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2617_ (.Y(_0784_),
    .A(\counter_lo_i.compare_value_i [15]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2618_ (.Y(_0785_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout18 (.X(net18),
    .A(net105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2620_ (.Y(_0787_),
    .B1(net50),
    .B2(\prescaler_lo_i.compare_value_i [7]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2621_ (.B(_0784_),
    .C(_0785_),
    .A(_0783_),
    .Y(_0788_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0787_));
 sg13g2_nor2b_2 _2622_ (.A(net23),
    .B_N(_0788_),
    .Y(r_rdata_o[15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2623_ (.Y(_0789_),
    .A(\prescaler_hi_i.compare_value_i [6]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2624_ (.Y(_0790_),
    .A(\counter_lo_i.compare_value_i [14]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2625_ (.Y(_0791_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2626_ (.Y(_0792_),
    .B1(net52),
    .B2(\prescaler_lo_i.compare_value_i [6]),
    .A2(net33),
    .A1(\counter_hi_i.compare_value_i [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2627_ (.B(_0790_),
    .C(_0791_),
    .A(_0789_),
    .Y(_0793_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0792_));
 sg13g2_nor2b_2 _2628_ (.A(net22),
    .B_N(_0793_),
    .Y(r_rdata_o[14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout17 (.A(_1020_),
    .X(net17),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout16 (.A(net105),
    .X(net16),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2631_ (.Y(_0796_),
    .A(\prescaler_hi_i.compare_value_i [5]),
    .B(net58),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2632_ (.Y(_0797_),
    .A(\counter_lo_i.compare_value_i [13]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout15 (.A(net105),
    .X(net15),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout14 (.A(net105),
    .X(net14),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2635_ (.Y(_0800_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout13 (.X(net13),
    .A(net105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2637_ (.Y(_0802_),
    .B1(net53),
    .B2(\prescaler_lo_i.compare_value_i [5]),
    .A2(net33),
    .A1(\counter_hi_i.compare_value_i [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2638_ (.B(_0797_),
    .C(_0800_),
    .A(_0796_),
    .Y(_0803_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0802_));
 sg13g2_nor2b_2 _2639_ (.A(net23),
    .B_N(_0803_),
    .Y(r_rdata_o[13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2640_ (.Y(_0804_),
    .A(\prescaler_hi_i.compare_value_i [4]),
    .B(net58),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout12 (.A(net105),
    .X(net12),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2642_ (.Y(_0806_),
    .A(\counter_lo_i.compare_value_i [12]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2643_ (.Y(_0807_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2644_ (.Y(_0808_),
    .B1(net53),
    .B2(\prescaler_lo_i.compare_value_i [4]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2645_ (.B(_0806_),
    .C(_0807_),
    .A(_0804_),
    .Y(_0809_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0808_));
 sg13g2_nor2b_2 _2646_ (.A(net23),
    .B_N(_0809_),
    .Y(r_rdata_o[12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2647_ (.Y(_0810_),
    .A(s_cfg_hi_reg[29]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2648_ (.Y(_0811_),
    .A(\counter_lo_i.compare_value_i [29]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2649_ (.Y(_0812_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2650_ (.Y(_0813_),
    .B1(net49),
    .B2(s_cfg_lo_reg[29]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2651_ (.B(_0811_),
    .C(_0812_),
    .A(_0810_),
    .Y(_0814_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0813_));
 sg13g2_nor2b_2 _2652_ (.A(net21),
    .B_N(_0814_),
    .Y(r_rdata_o[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2653_ (.Y(_0815_),
    .A(\prescaler_hi_i.compare_value_i [3]),
    .B(net58),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2654_ (.Y(_0816_),
    .A(\counter_lo_i.compare_value_i [11]),
    .B(net38),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2655_ (.Y(_0817_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2656_ (.Y(_0818_),
    .B1(net52),
    .B2(\prescaler_lo_i.compare_value_i [3]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2657_ (.B(_0816_),
    .C(_0817_),
    .A(_0815_),
    .Y(_0819_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0818_));
 sg13g2_nor2b_2 _2658_ (.A(net24),
    .B_N(_0819_),
    .Y(r_rdata_o[11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2659_ (.Y(_0820_),
    .A(\prescaler_hi_i.compare_value_i [2]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2660_ (.Y(_0821_),
    .A(\counter_lo_i.compare_value_i [10]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2661_ (.Y(_0822_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2662_ (.Y(_0823_),
    .B1(net52),
    .B2(\prescaler_lo_i.compare_value_i [2]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2663_ (.B(_0821_),
    .C(_0822_),
    .A(_0820_),
    .Y(_0824_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0823_));
 sg13g2_nor2b_2 _2664_ (.A(net24),
    .B_N(_0824_),
    .Y(r_rdata_o[10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2665_ (.Y(_0825_),
    .A(\prescaler_hi_i.compare_value_i [1]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2666_ (.Y(_0826_),
    .A(\counter_lo_i.compare_value_i [9]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2667_ (.Y(_0827_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2668_ (.Y(_0828_),
    .B1(net52),
    .B2(\prescaler_lo_i.compare_value_i [1]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2669_ (.B(_0826_),
    .C(_0827_),
    .A(_0825_),
    .Y(_0829_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0828_));
 sg13g2_nor2b_2 _2670_ (.A(net23),
    .B_N(_0829_),
    .Y(r_rdata_o[9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2671_ (.Y(_0830_),
    .A(\prescaler_hi_i.compare_value_i [0]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2672_ (.Y(_0831_),
    .A(\counter_lo_i.compare_value_i [8]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2673_ (.Y(_0832_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2674_ (.Y(_0833_),
    .B1(net52),
    .B2(\prescaler_lo_i.compare_value_i [0]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2675_ (.B(_0831_),
    .C(_0832_),
    .A(_0830_),
    .Y(_0834_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0833_));
 sg13g2_nor2b_2 _2676_ (.A(net22),
    .B_N(_0834_),
    .Y(r_rdata_o[8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2677_ (.Y(_0835_),
    .A(s_cfg_hi_reg[7]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2678_ (.Y(_0836_),
    .A(\counter_lo_i.compare_value_i [7]),
    .B(net36),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2679_ (.Y(_0837_),
    .B1(net42),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .A2(net47),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2680_ (.Y(_0838_),
    .B1(net52),
    .B2(s_cfg_lo_reg[7]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2681_ (.B(_0836_),
    .C(_0837_),
    .A(_0835_),
    .Y(_0839_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0838_));
 sg13g2_nor2b_2 _2682_ (.A(net24),
    .B_N(_0839_),
    .Y(r_rdata_o[7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2683_ (.Y(_0840_),
    .A(s_cfg_hi_reg[6]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2684_ (.Y(_0841_),
    .A(\counter_lo_i.compare_value_i [6]),
    .B(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2685_ (.Y(_0842_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout11 (.A(net105),
    .X(net11),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2687_ (.Y(_0844_),
    .B1(net51),
    .B2(s_cfg_lo_reg[6]),
    .A2(net32),
    .A1(\counter_hi_i.compare_value_i [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2688_ (.B(_0841_),
    .C(_0842_),
    .A(_0840_),
    .Y(_0845_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0844_));
 sg13g2_nor2b_2 _2689_ (.A(net24),
    .B_N(_0845_),
    .Y(r_rdata_o[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2690_ (.Y(_0846_),
    .A(s_cfg_hi_reg[5]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2691_ (.Y(_0847_),
    .A(\counter_lo_i.compare_value_i [5]),
    .B(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2692_ (.Y(_0848_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2693_ (.Y(_0849_),
    .B1(net51),
    .B2(s_cfg_lo_reg[5]),
    .A2(net31),
    .A1(\counter_hi_i.compare_value_i [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2694_ (.B(_0847_),
    .C(_0848_),
    .A(_0846_),
    .Y(_0850_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0849_));
 sg13g2_nor2b_2 _2695_ (.A(net23),
    .B_N(_0850_),
    .Y(r_rdata_o[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout10 (.A(net105),
    .X(net10),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2697_ (.Y(_0852_),
    .A(\counter_hi_i.compare_value_i [4]),
    .B(net31),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2698_ (.Y(_0853_),
    .A(\counter_lo_i.compare_value_i [4]),
    .B(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout9 (.A(_0960_),
    .X(net9),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout8 (.A(_0960_),
    .X(net8),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2701_ (.Y(_0856_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout7 (.A(_0960_),
    .X(net7),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2703_ (.Y(_0858_),
    .B1(net52),
    .B2(s_cfg_lo_reg[4]),
    .A2(net56),
    .A1(s_cfg_hi_reg[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2704_ (.B(_0853_),
    .C(_0856_),
    .A(_0852_),
    .Y(_0859_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0858_));
 sg13g2_nor2b_2 _2705_ (.A(net25),
    .B_N(_0859_),
    .Y(r_rdata_o[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout6 (.A(_0960_),
    .X(net6),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2707_ (.Y(_0861_),
    .A(s_cfg_hi_reg[3]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout5 (.A(_0260_),
    .X(net5),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2709_ (.Y(_0863_),
    .A(\counter_lo_i.compare_value_i [3]),
    .B(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2710_ (.Y(_0864_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2711_ (.Y(_0865_),
    .B1(net51),
    .B2(s_cfg_lo_reg[3]),
    .A2(net31),
    .A1(\counter_hi_i.compare_value_i [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2712_ (.B(_0863_),
    .C(_0864_),
    .A(_0861_),
    .Y(_0866_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0865_));
 sg13g2_nor2b_2 _2713_ (.A(net22),
    .B_N(_0866_),
    .Y(r_rdata_o[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2714_ (.Y(_0867_),
    .A(s_cfg_hi_reg[2]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2715_ (.Y(_0868_),
    .A(\counter_lo_i.compare_value_i [2]),
    .B(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2716_ (.Y(_0869_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2717_ (.Y(_0870_),
    .B1(net51),
    .B2(s_cfg_lo_reg[2]),
    .A2(net31),
    .A1(\counter_hi_i.compare_value_i [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2718_ (.B(_0868_),
    .C(_0869_),
    .A(_0867_),
    .Y(_0871_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0870_));
 sg13g2_nor2b_2 _2719_ (.A(net24),
    .B_N(_0871_),
    .Y(r_rdata_o[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2720_ (.Y(_0872_),
    .A(s_cfg_hi_reg[28]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2721_ (.Y(_0873_),
    .A(\counter_lo_i.compare_value_i [28]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2722_ (.Y(_0874_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2723_ (.Y(_0875_),
    .B1(net49),
    .B2(s_cfg_lo_reg[28]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2724_ (.B(_0873_),
    .C(_0874_),
    .A(_0872_),
    .Y(_0876_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0875_));
 sg13g2_nor2b_2 _2725_ (.A(net21),
    .B_N(_0876_),
    .Y(r_rdata_o[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2726_ (.Y(_0877_),
    .A(s_cfg_hi_reg[1]),
    .B(net57),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2727_ (.Y(_0878_),
    .A(\counter_lo_i.compare_value_i [1]),
    .B(net37),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2728_ (.Y(_0879_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2729_ (.Y(_0880_),
    .B1(net51),
    .B2(s_cfg_lo_reg[1]),
    .A2(net31),
    .A1(\counter_hi_i.compare_value_i [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2730_ (.B(_0878_),
    .C(_0879_),
    .A(_0877_),
    .Y(_0881_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0880_));
 sg13g2_nor2b_2 _2731_ (.A(net25),
    .B_N(_0881_),
    .Y(r_rdata_o[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2732_ (.Y(_0882_),
    .A(s_cfg_hi_reg[0]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2733_ (.Y(_0883_),
    .A(\counter_hi_i.compare_value_i [0]),
    .B(net31),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2734_ (.Y(_0884_),
    .B1(net41),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .A2(net46),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2735_ (.Y(_0885_),
    .B1(net51),
    .B2(s_cfg_lo_reg[0]),
    .A2(net37),
    .A1(\counter_lo_i.compare_value_i [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2736_ (.B(_0883_),
    .C(_0884_),
    .A(_0882_),
    .Y(_0886_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0885_));
 sg13g2_nor2b_2 _2737_ (.A(net23),
    .B_N(_0886_),
    .Y(r_rdata_o[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2738_ (.Y(_0887_),
    .A(s_cfg_hi_reg[27]),
    .B(net56),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2739_ (.Y(_0888_),
    .A(\counter_lo_i.compare_value_i [27]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2740_ (.Y(_0889_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2741_ (.Y(_0890_),
    .B1(net49),
    .B2(s_cfg_lo_reg[27]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2742_ (.B(_0888_),
    .C(_0889_),
    .A(_0887_),
    .Y(_0891_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0890_));
 sg13g2_nor2b_2 _2743_ (.A(net22),
    .B_N(_0891_),
    .Y(r_rdata_o[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2744_ (.Y(_0892_),
    .A(s_cfg_hi_reg[26]),
    .B(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2745_ (.Y(_0893_),
    .A(\counter_lo_i.compare_value_i [26]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2746_ (.Y(_0894_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2747_ (.Y(_0895_),
    .B1(net50),
    .B2(s_cfg_lo_reg[26]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2748_ (.B(_0893_),
    .C(_0894_),
    .A(_0892_),
    .Y(_0896_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0895_));
 sg13g2_nor2b_2 _2749_ (.A(net24),
    .B_N(_0896_),
    .Y(r_rdata_o[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2750_ (.Y(_0897_),
    .A(s_cfg_hi_reg[25]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2751_ (.Y(_0898_),
    .A(\counter_lo_i.compare_value_i [25]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2752_ (.Y(_0899_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2753_ (.Y(_0900_),
    .B1(net49),
    .B2(s_cfg_lo_reg[25]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2754_ (.B(_0898_),
    .C(_0899_),
    .A(_0897_),
    .Y(_0901_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0900_));
 sg13g2_nor2b_2 _2755_ (.A(net24),
    .B_N(_0901_),
    .Y(r_rdata_o[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2756_ (.Y(_0902_),
    .A(s_cfg_hi_reg[24]),
    .B(net55),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2757_ (.Y(_0903_),
    .A(\counter_lo_i.compare_value_i [24]),
    .B(net35),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2758_ (.Y(_0904_),
    .B1(net40),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .A2(net45),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2759_ (.Y(_0905_),
    .B1(net50),
    .B2(s_cfg_lo_reg[24]),
    .A2(net30),
    .A1(\counter_hi_i.compare_value_i [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2760_ (.B(_0903_),
    .C(_0904_),
    .A(_0902_),
    .Y(_0906_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0905_));
 sg13g2_nor2b_2 _2761_ (.A(net21),
    .B_N(_0906_),
    .Y(r_rdata_o[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2762_ (.Y(_0907_),
    .A(s_cfg_hi_reg[23]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2763_ (.Y(_0908_),
    .A(\counter_lo_i.compare_value_i [23]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2764_ (.Y(_0909_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2765_ (.Y(_0910_),
    .B1(net49),
    .B2(s_cfg_lo_reg[23]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2766_ (.B(_0908_),
    .C(_0909_),
    .A(_0907_),
    .Y(_0911_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0910_));
 sg13g2_nor2b_2 _2767_ (.A(net21),
    .B_N(_0911_),
    .Y(r_rdata_o[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2768_ (.Y(_0912_),
    .A(s_cfg_hi_reg[22]),
    .B(net54),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2769_ (.Y(_0913_),
    .A(\counter_lo_i.compare_value_i [22]),
    .B(net34),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2770_ (.Y(_0914_),
    .B1(net39),
    .B2(\counter_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .A2(net44),
    .A1(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2771_ (.Y(_0915_),
    .B1(net49),
    .B2(s_cfg_lo_reg[22]),
    .A2(net29),
    .A1(\counter_hi_i.compare_value_i [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _2772_ (.B(_0913_),
    .C(_0914_),
    .A(_0912_),
    .Y(_0916_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_0915_));
 sg13g2_nor2b_2 _2773_ (.A(net21),
    .B_N(_0916_),
    .Y(r_rdata_o[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2774_ (.A0(wdata_i[5]),
    .A1(s_cfg_hi_reg[5]),
    .S(net90),
    .X(s_cfg_hi[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 _2775_ (.VDD(VDD),
    .Y(_0917_),
    .A(\counter_hi_i.target_reached_o ),
    .VSS(VSS));
 sg13g2_mux2_1 _2776_ (.A0(s_cfg_lo_reg[5]),
    .A1(wdata_i[5]),
    .S(net84),
    .X(s_cfg_lo[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a22oi_1 _2777_ (.Y(_0918_),
    .B1(s_cfg_lo[5]),
    .B2(\counter_lo_i.target_reached_o ),
    .A2(s_cfg_hi[5]),
    .A1(\s_cfg_hi_$_OR__Y_A_$_MUX__Y_S_$_AND__Y_A_$_AND__Y_A ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2778_ (.A0(wdata_i[0]),
    .A1(s_cfg_hi_reg[0]),
    .S(net90),
    .X(_0919_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2779_ (.B1(_0919_),
    .VDD(VDD),
    .Y(_0920_),
    .VSS(VSS),
    .A1(_0917_),
    .A2(_0918_));
 sg13g2_a22oi_1 _2780_ (.Y(_0921_),
    .B1(s_cfg_hi[3]),
    .B2(event_hi_i),
    .A2(_1141_),
    .A1(_0938_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2781_ (.Y(s_cfg_hi[0]),
    .A(_0920_),
    .B(_0921_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2782_ (.A0(wdata_i[16]),
    .A1(s_cfg_hi_reg[16]),
    .S(net90),
    .X(_0080_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2783_ (.A0(wdata_i[17]),
    .A1(s_cfg_hi_reg[17]),
    .S(net89),
    .X(_0081_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2784_ (.A0(wdata_i[18]),
    .A1(s_cfg_hi_reg[18]),
    .S(net89),
    .X(_0082_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2785_ (.A0(wdata_i[19]),
    .A1(s_cfg_hi_reg[19]),
    .S(net89),
    .X(_0083_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _2786_ (.A(_0233_),
    .B(net75),
    .C(net90),
    .Y(_0084_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2787_ (.A0(wdata_i[20]),
    .A1(s_cfg_hi_reg[20]),
    .S(net89),
    .X(_0085_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2788_ (.A0(wdata_i[21]),
    .A1(s_cfg_hi_reg[21]),
    .S(net88),
    .X(_0086_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2789_ (.A0(wdata_i[22]),
    .A1(s_cfg_hi_reg[22]),
    .S(net88),
    .X(_0087_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2790_ (.A0(wdata_i[23]),
    .A1(s_cfg_hi_reg[23]),
    .S(net88),
    .X(_0088_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2791_ (.A0(wdata_i[24]),
    .A1(s_cfg_hi_reg[24]),
    .S(net89),
    .X(_0089_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout4 (.A(_1172_),
    .X(net4),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2793_ (.A0(wdata_i[25]),
    .A1(s_cfg_hi_reg[25]),
    .S(net88),
    .X(_0090_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2794_ (.Y(_0923_),
    .A(s_cfg_hi_reg[26]),
    .B(net89),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2795_ (.B1(_0923_),
    .VDD(VDD),
    .Y(_0091_),
    .VSS(VSS),
    .A1(_1153_),
    .A2(net89));
 sg13g2_mux2_1 _2796_ (.A0(wdata_i[27]),
    .A1(s_cfg_hi_reg[27]),
    .S(net88),
    .X(_0092_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2797_ (.A0(wdata_i[28]),
    .A1(s_cfg_hi_reg[28]),
    .S(net88),
    .X(_0093_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2798_ (.A0(wdata_i[29]),
    .A1(s_cfg_hi_reg[29]),
    .S(net88),
    .X(_0094_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2799_ (.A0(wdata_i[2]),
    .A1(s_cfg_hi_reg[2]),
    .S(net91),
    .X(_0095_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2800_ (.A0(wdata_i[30]),
    .A1(s_cfg_hi_reg[30]),
    .S(net88),
    .X(_0096_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2801_ (.A0(wdata_i[31]),
    .A1(s_cfg_hi_reg[31]),
    .S(net90),
    .X(_0097_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2802_ (.A0(wdata_i[4]),
    .A1(s_cfg_hi_reg[4]),
    .S(net90),
    .X(_0098_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2803_ (.A0(wdata_i[6]),
    .A1(s_cfg_hi_reg[6]),
    .S(net90),
    .X(_0099_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2804_ (.A0(wdata_i[7]),
    .A1(s_cfg_hi_reg[7]),
    .S(net92),
    .X(_0100_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2b_1 _2805_ (.A(_0239_),
    .B_N(s_cfg_lo[5]),
    .Y(_0924_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2806_ (.A(_0935_),
    .B(net85),
    .Y(_0925_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _2807_ (.VSS(VSS),
    .VDD(VDD),
    .A1(wdata_i[0]),
    .A2(net85),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_a22oi_1 _2808_ (.Y(_0927_),
    .B1(s_cfg_lo[3]),
    .B2(event_lo_i),
    .A2(_0246_),
    .A1(_0938_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2809_ (.B1(_0927_),
    .VDD(VDD),
    .Y(s_cfg_lo[0]),
    .VSS(VSS),
    .A1(_0924_),
    .A2(_0926_));
 sg13g2_mux2_1 _2810_ (.A0(s_cfg_lo_reg[16]),
    .A1(wdata_i[16]),
    .S(net84),
    .X(_0101_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2811_ (.A0(s_cfg_lo_reg[17]),
    .A1(wdata_i[17]),
    .S(net83),
    .X(_0102_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout3 (.A(_1172_),
    .X(net3),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2813_ (.A0(s_cfg_lo_reg[18]),
    .A1(wdata_i[18]),
    .S(net83),
    .X(_0103_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2814_ (.A0(s_cfg_lo_reg[19]),
    .A1(wdata_i[19]),
    .S(net83),
    .X(_0104_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2815_ (.Y(_0929_),
    .A(wdata_i[1]),
    .B(net85),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _2816_ (.A(net73),
    .B(_0929_),
    .Y(_0105_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2817_ (.A0(s_cfg_lo_reg[20]),
    .A1(wdata_i[20]),
    .S(net83),
    .X(_0106_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2818_ (.A0(s_cfg_lo_reg[21]),
    .A1(wdata_i[21]),
    .S(net82),
    .X(_0107_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2819_ (.A0(s_cfg_lo_reg[22]),
    .A1(wdata_i[22]),
    .S(net82),
    .X(_0108_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2820_ (.A0(s_cfg_lo_reg[23]),
    .A1(wdata_i[23]),
    .S(net82),
    .X(_0109_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2821_ (.A0(s_cfg_lo_reg[24]),
    .A1(wdata_i[24]),
    .S(net83),
    .X(_0110_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2822_ (.A0(s_cfg_lo_reg[25]),
    .A1(wdata_i[25]),
    .S(net82),
    .X(_0111_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2823_ (.A0(s_cfg_lo_reg[26]),
    .A1(wdata_i[26]),
    .S(net83),
    .X(_0112_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2824_ (.A0(s_cfg_lo_reg[27]),
    .A1(wdata_i[27]),
    .S(net82),
    .X(_0113_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2825_ (.A0(s_cfg_lo_reg[28]),
    .A1(wdata_i[28]),
    .S(net82),
    .X(_0114_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_mux2_1 _2826_ (.A0(s_cfg_lo_reg[29]),
    .A1(wdata_i[29]),
    .S(net82),
    .X(_0115_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2827_ (.Y(_0930_),
    .A(wdata_i[2]),
    .B(net84),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2828_ (.B1(_0930_),
    .VDD(VDD),
    .Y(_0116_),
    .VSS(VSS),
    .A1(_0470_),
    .A2(net84));
 sg13g2_mux2_1 _2829_ (.A0(s_cfg_lo_reg[30]),
    .A1(wdata_i[30]),
    .S(net82),
    .X(_0117_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2830_ (.Y(_0931_),
    .A(wdata_i[31]),
    .B(net84),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2831_ (.B1(_0931_),
    .VDD(VDD),
    .Y(_0118_),
    .VSS(VSS),
    .A1(_0238_),
    .A2(net84));
 sg13g2_nand2_1 _2832_ (.Y(_0932_),
    .A(wdata_i[4]),
    .B(net85),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2833_ (.B1(_0932_),
    .VDD(VDD),
    .Y(_0119_),
    .VSS(VSS),
    .A1(_0237_),
    .A2(net85));
 sg13g2_mux2_1 _2834_ (.A0(s_cfg_lo_reg[6]),
    .A1(wdata_i[6]),
    .S(net84),
    .X(_0120_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2_1 _2835_ (.Y(_0933_),
    .A(wdata_i[7]),
    .B(net86),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _2836_ (.B1(_0933_),
    .VDD(VDD),
    .Y(_0121_),
    .VSS(VSS),
    .A1(_0985_),
    .A2(net86));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net91),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tiehi timer_unit_2 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net2));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[0]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0000_),
    .Q_N(_1334_),
    .Q(\counter_hi_i.compare_value_i [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[10]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0001_),
    .Q_N(_1333_),
    .Q(\counter_hi_i.compare_value_i [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[11]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0002_),
    .Q_N(_1332_),
    .Q(\counter_hi_i.compare_value_i [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[12]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0003_),
    .Q(\counter_hi_i.compare_value_i [12]),
    .Q_N(_1331_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[13]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0004_),
    .Q(\counter_hi_i.compare_value_i [13]),
    .Q_N(_1330_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[14]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0005_),
    .Q(\counter_hi_i.compare_value_i [14]),
    .Q_N(_1329_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[15]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0006_),
    .Q_N(_1328_),
    .Q(\counter_hi_i.compare_value_i [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[16]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(_0007_),
    .Q_N(_1327_),
    .Q(\counter_hi_i.compare_value_i [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[17]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0008_),
    .Q(\counter_hi_i.compare_value_i [17]),
    .Q_N(_1326_),
    .CLK(clknet_leaf_36_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[18]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0009_),
    .Q_N(_1325_),
    .Q(\counter_hi_i.compare_value_i [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[19]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0010_),
    .Q_N(_1324_),
    .Q(\counter_hi_i.compare_value_i [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[1]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0011_),
    .Q_N(_1323_),
    .Q(\counter_hi_i.compare_value_i [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[20]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0012_),
    .Q_N(_1322_),
    .Q(\counter_hi_i.compare_value_i [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[21]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0013_),
    .Q(\counter_hi_i.compare_value_i [21]),
    .Q_N(_1321_),
    .CLK(clknet_leaf_27_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[22]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0014_),
    .Q(\counter_hi_i.compare_value_i [22]),
    .Q_N(_1320_),
    .CLK(clknet_leaf_28_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[23]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0015_),
    .Q_N(_1319_),
    .Q(\counter_hi_i.compare_value_i [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[24]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0016_),
    .Q(\counter_hi_i.compare_value_i [24]),
    .Q_N(_1318_),
    .CLK(clknet_leaf_29_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[25]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0017_),
    .Q(\counter_hi_i.compare_value_i [25]),
    .Q_N(_1317_),
    .CLK(clknet_leaf_29_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[26]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0018_),
    .Q(\counter_hi_i.compare_value_i [26]),
    .Q_N(_1316_),
    .CLK(clknet_leaf_29_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[27]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0019_),
    .Q_N(_1315_),
    .Q(\counter_hi_i.compare_value_i [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[28]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0020_),
    .Q_N(_1314_),
    .Q(\counter_hi_i.compare_value_i [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[29]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0021_),
    .Q_N(_1313_),
    .Q(\counter_hi_i.compare_value_i [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[2]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0022_),
    .Q_N(_1312_),
    .Q(\counter_hi_i.compare_value_i [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[30]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0023_),
    .Q_N(_1311_),
    .Q(\counter_hi_i.compare_value_i [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[31]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0024_),
    .Q_N(_1310_),
    .Q(\counter_hi_i.compare_value_i [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[3]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0025_),
    .Q_N(_1309_),
    .Q(\counter_hi_i.compare_value_i [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[4]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(_0026_),
    .Q_N(_1308_),
    .Q(\counter_hi_i.compare_value_i [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[5]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0027_),
    .Q_N(_1307_),
    .Q(\counter_hi_i.compare_value_i [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[6]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(_0028_),
    .Q_N(_1306_),
    .Q(\counter_hi_i.compare_value_i [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[7]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0029_),
    .Q_N(_1305_),
    .Q(\counter_hi_i.compare_value_i [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.compare_value_i[8]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(_0030_),
    .Q_N(_1304_),
    .Q(\counter_hi_i.compare_value_i [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.compare_value_i[9]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0031_),
    .Q(\counter_hi_i.compare_value_i [9]),
    .Q_N(_1335_),
    .CLK(clknet_leaf_3_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [0]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__S_31_B [0]),
    .CLK(clknet_leaf_1_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[10]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [10]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .Q_N(_1336_),
    .CLK(clknet_leaf_3_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[11]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [11]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .Q_N(_1337_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[12]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [12]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .Q_N(_1338_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[13]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [13]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .Q_N(_1339_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[14]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [14]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .Q_N(_1340_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[15]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [15]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .Q_N(_1341_),
    .CLK(clknet_leaf_35_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[16]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [16]),
    .Q_N(_1342_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[17]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [17]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .Q_N(_1343_),
    .CLK(clknet_leaf_35_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[18]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [18]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .Q_N(_1344_),
    .CLK(clknet_leaf_32_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[19]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [19]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .Q_N(_1345_),
    .CLK(clknet_leaf_32_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[1]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [1]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .Q_N(_1346_),
    .CLK(clknet_leaf_38_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[20]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [20]),
    .Q_N(_1347_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[21]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [21]),
    .Q_N(_1348_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[22]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [22]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .Q_N(_1349_),
    .CLK(clknet_leaf_25_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[23]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [23]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .Q_N(_1350_),
    .CLK(clknet_leaf_28_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[24]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [24]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .Q_N(_1351_),
    .CLK(clknet_leaf_28_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[25]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [25]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .Q_N(_1352_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[26]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [26]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .Q_N(_1353_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[27]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [27]),
    .Q_N(_1354_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[28]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [28]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .Q_N(_1355_),
    .CLK(clknet_leaf_27_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[29]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [29]),
    .Q_N(_1356_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[2]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [2]),
    .Q_N(_1357_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[30]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [30]),
    .Q_N(_1358_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[31]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [31]),
    .Q_N(_1359_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[3]_reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [3]),
    .Q_N(_1360_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[4]_reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [4]),
    .Q_N(_1361_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[5]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [5]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .Q_N(_1362_),
    .CLK(clknet_leaf_38_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[6]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [6]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .Q_N(_1363_),
    .CLK(clknet_leaf_37_clk_i));
 sg13g2_dfrbp_2 \counter_hi_i.counter_value_o[7]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_hi_i.s_count [7]),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .Q_N(_1364_),
    .CLK(clknet_leaf_36_clk_i));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[8]_reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [8]),
    .Q_N(_1365_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.counter_value_o[9]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.s_count [9]),
    .Q_N(_1366_),
    .Q(\counter_hi_i.enable_count_i_$_MUX__S_31_B [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_hi_i.target_reached_o_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_hi_i.target_reached_o_reg_D ),
    .Q_N(_1303_),
    .Q(\counter_hi_i.target_reached_o ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[0]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0032_),
    .Q_N(_1302_),
    .Q(\counter_lo_i.compare_value_i [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[10]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0033_),
    .Q_N(_1301_),
    .Q(\counter_lo_i.compare_value_i [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[11]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0034_),
    .Q_N(_1300_),
    .Q(\counter_lo_i.compare_value_i [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[12]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0035_),
    .Q_N(_1299_),
    .Q(\counter_lo_i.compare_value_i [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[13]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0036_),
    .Q_N(_1298_),
    .Q(\counter_lo_i.compare_value_i [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[14]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(_0037_),
    .Q_N(_1297_),
    .Q(\counter_lo_i.compare_value_i [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[15]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0038_),
    .Q_N(_1296_),
    .Q(\counter_lo_i.compare_value_i [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[16]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(_0039_),
    .Q_N(_1295_),
    .Q(\counter_lo_i.compare_value_i [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[17]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0040_),
    .Q_N(_1294_),
    .Q(\counter_lo_i.compare_value_i [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[18]_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(rst_ni),
    .D(_0041_),
    .Q_N(_1293_),
    .Q(\counter_lo_i.compare_value_i [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[19]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0042_),
    .Q_N(_1292_),
    .Q(\counter_lo_i.compare_value_i [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[1]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0043_),
    .Q_N(_1291_),
    .Q(\counter_lo_i.compare_value_i [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[20]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0044_),
    .Q_N(_1290_),
    .Q(\counter_lo_i.compare_value_i [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[21]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0045_),
    .Q_N(_1289_),
    .Q(\counter_lo_i.compare_value_i [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[22]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0046_),
    .Q_N(_1288_),
    .Q(\counter_lo_i.compare_value_i [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[23]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0047_),
    .Q_N(_1287_),
    .Q(\counter_lo_i.compare_value_i [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[24]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0048_),
    .Q_N(_1286_),
    .Q(\counter_lo_i.compare_value_i [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[25]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0049_),
    .Q_N(_1285_),
    .Q(\counter_lo_i.compare_value_i [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[26]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0050_),
    .Q_N(_1284_),
    .Q(\counter_lo_i.compare_value_i [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[27]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0051_),
    .Q_N(_1283_),
    .Q(\counter_lo_i.compare_value_i [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[28]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(_0052_),
    .Q_N(_1282_),
    .Q(\counter_lo_i.compare_value_i [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[29]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0053_),
    .Q_N(_1281_),
    .Q(\counter_lo_i.compare_value_i [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[2]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0054_),
    .Q_N(_1280_),
    .Q(\counter_lo_i.compare_value_i [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[30]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0055_),
    .Q_N(_1279_),
    .Q(\counter_lo_i.compare_value_i [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[31]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(_0056_),
    .Q_N(_1278_),
    .Q(\counter_lo_i.compare_value_i [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[3]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0057_),
    .Q_N(_1277_),
    .Q(\counter_lo_i.compare_value_i [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[4]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0058_),
    .Q_N(_1276_),
    .Q(\counter_lo_i.compare_value_i [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[5]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0059_),
    .Q_N(_1275_),
    .Q(\counter_lo_i.compare_value_i [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[6]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(_0060_),
    .Q_N(_1274_),
    .Q(\counter_lo_i.compare_value_i [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[7]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0061_),
    .Q_N(_1273_),
    .Q(\counter_lo_i.compare_value_i [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.compare_value_i[8]_reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(rst_ni),
    .D(_0062_),
    .Q_N(_1272_),
    .Q(\counter_lo_i.compare_value_i [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.compare_value_i[9]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0063_),
    .Q(\counter_lo_i.compare_value_i [9]),
    .Q_N(_1367_),
    .CLK(clknet_leaf_13_clk_i));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [0]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_A ),
    .CLK(clknet_leaf_7_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[10]_reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [10]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_10_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[11]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [11]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_10_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[12]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [12]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_9_A ),
    .CLK(clknet_leaf_4_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[13]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [13]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_9_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[14]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [14]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_8_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[15]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [15]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_8_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[16]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [16]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_7_A ),
    .CLK(clknet_leaf_4_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[17]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [17]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_7_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[18]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [18]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_6_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[19]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [19]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_6_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[1]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [1]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_15_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[20]_reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [20]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_5_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[21]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [21]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_5_B ),
    .CLK(clknet_leaf_25_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[22]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [22]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_4_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[23]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [23]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_4_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[24]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [24]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_3_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[25]_reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [25]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_3_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[26]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [26]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_2_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[27]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [27]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_2_B ),
    .CLK(clknet_leaf_23_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[28]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [28]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_1_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[29]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [29]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_1_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[2]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [2]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_14_A ),
    .CLK(clknet_leaf_7_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[30]_reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [30]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[31]_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [31]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[3]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [3]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_14_B ),
    .CLK(clknet_leaf_8_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[4]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [4]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_13_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[5]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [5]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_13_B ),
    .CLK(clknet_leaf_6_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.counter_value_o[6]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.s_count [6]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_12_A ),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[7]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [7]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_12_B ),
    .CLK(clknet_leaf_4_clk_i));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[8]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [8]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_11_A ),
    .CLK(clknet_leaf_5_clk_i));
 sg13g2_dfrbp_2 \counter_lo_i.counter_value_o[9]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\counter_lo_i.s_count [9]),
    .Q(\counter_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .Q_N(\counter_hi_i.enable_count_i_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_11_B ),
    .CLK(clknet_leaf_5_clk_i));
 sg13g2_dfrbp_1 \counter_lo_i.target_reached_o_reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(rst_ni),
    .D(\counter_lo_i.target_reached_o_reg_D ),
    .Q_N(_1271_),
    .Q(\counter_lo_i.target_reached_o ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.compare_value_i[0]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0064_),
    .Q_N(_1270_),
    .Q(\prescaler_hi_i.compare_value_i [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.compare_value_i[1]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0065_),
    .Q_N(_1269_),
    .Q(\prescaler_hi_i.compare_value_i [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.compare_value_i[2]_reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(rst_ni),
    .D(_0066_),
    .Q_N(_1268_),
    .Q(\prescaler_hi_i.compare_value_i [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.compare_value_i[3]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0067_),
    .Q_N(_1267_),
    .Q(\prescaler_hi_i.compare_value_i [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.compare_value_i[4]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0068_),
    .Q_N(_1266_),
    .Q(\prescaler_hi_i.compare_value_i [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_hi_i.compare_value_i[5]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0069_),
    .Q(\prescaler_hi_i.compare_value_i [5]),
    .Q_N(_1265_),
    .CLK(clknet_leaf_16_clk_i));
 sg13g2_dfrbp_2 \prescaler_hi_i.compare_value_i[6]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0070_),
    .Q(\prescaler_hi_i.compare_value_i [6]),
    .Q_N(_1264_),
    .CLK(clknet_leaf_15_clk_i));
 sg13g2_dfrbp_2 \prescaler_hi_i.compare_value_i[7]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0071_),
    .Q(\prescaler_hi_i.compare_value_i [7]),
    .Q_N(_1368_),
    .CLK(clknet_leaf_24_clk_i));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[0]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [0]),
    .Q_N(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [0]),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[10]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [10]),
    .Q_N(_1369_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_hi_i.counter_value_o[11]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_hi_i.s_count [11]),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [11]),
    .Q_N(_1370_),
    .CLK(clknet_leaf_21_clk_i));
 sg13g2_dfrbp_2 \prescaler_hi_i.counter_value_o[12]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_hi_i.s_count [12]),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [12]),
    .Q_N(_1371_),
    .CLK(clknet_leaf_18_clk_i));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[13]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [13]),
    .Q_N(_1372_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[14]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [14]),
    .Q_N(_1373_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[15]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [15]),
    .Q_N(_1374_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[16]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [16]),
    .Q_N(_1375_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[17]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [17]),
    .Q_N(_1376_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[18]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [18]),
    .Q_N(_1377_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[19]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [19]),
    .Q_N(_1378_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[1]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [1]),
    .Q_N(_1379_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[20]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [20]),
    .Q_N(_1380_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[21]_reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [21]),
    .Q_N(_1381_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_hi_i.counter_value_o[22]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_hi_i.s_count [22]),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [22]),
    .Q_N(_1382_),
    .CLK(clknet_leaf_20_clk_i));
 sg13g2_dfrbp_2 \prescaler_hi_i.counter_value_o[23]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_hi_i.s_count [23]),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [23]),
    .Q_N(_1383_),
    .CLK(clknet_leaf_20_clk_i));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[24]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [24]),
    .Q_N(_1384_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[25]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [25]),
    .Q_N(_1385_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[26]_reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [26]),
    .Q_N(_1386_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[27]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [27]),
    .Q_N(_1387_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[28]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [28]),
    .Q_N(_1388_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_hi_i.counter_value_o[29]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_hi_i.s_count [29]),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [29]),
    .Q_N(_1389_),
    .CLK(clknet_leaf_22_clk_i));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[2]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [2]),
    .Q_N(_1390_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[30]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [30]),
    .Q_N(_1391_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[31]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [31]),
    .Q_N(_1392_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[3]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [3]),
    .Q_N(_1393_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[4]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [4]),
    .Q_N(_1394_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[5]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [5]),
    .Q_N(_1395_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[6]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [6]),
    .Q_N(_1396_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[7]_reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [7]),
    .Q_N(_1397_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[8]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [8]),
    .Q_N(_1398_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [8]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.counter_value_o[9]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.s_count [9]),
    .Q_N(_1399_),
    .Q(\prescaler_hi_i.enable_count_i_$_MUX__S_31_B [9]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_hi_i.target_reached_o_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_hi_i.target_reached_o_reg_D ),
    .Q_N(_1263_),
    .Q(\prescaler_hi_i.target_reached_o ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.compare_value_i[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0072_),
    .Q(\prescaler_lo_i.compare_value_i [0]),
    .Q_N(_1262_),
    .CLK(clknet_leaf_10_clk_i));
 sg13g2_dfrbp_2 \prescaler_lo_i.compare_value_i[1]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0073_),
    .Q(\prescaler_lo_i.compare_value_i [1]),
    .Q_N(_1261_),
    .CLK(clknet_leaf_11_clk_i));
 sg13g2_dfrbp_2 \prescaler_lo_i.compare_value_i[2]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0074_),
    .Q(\prescaler_lo_i.compare_value_i [2]),
    .Q_N(_1260_),
    .CLK(clknet_leaf_13_clk_i));
 sg13g2_dfrbp_2 \prescaler_lo_i.compare_value_i[3]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0075_),
    .Q(\prescaler_lo_i.compare_value_i [3]),
    .Q_N(_1259_),
    .CLK(clknet_leaf_13_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.compare_value_i[4]_reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(rst_ni),
    .D(_0076_),
    .Q_N(_1258_),
    .Q(\prescaler_lo_i.compare_value_i [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.compare_value_i[5]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0077_),
    .Q_N(_1257_),
    .Q(\prescaler_lo_i.compare_value_i [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.compare_value_i[6]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(_0078_),
    .Q_N(_1256_),
    .Q(\prescaler_lo_i.compare_value_i [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.compare_value_i[7]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0079_),
    .Q_N(_1400_),
    .Q(\prescaler_lo_i.compare_value_i [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[0]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [0]),
    .Q_N(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [0]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_B_$_XOR__Y_B [0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[10]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [10]),
    .Q_N(_1401_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [10]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[11]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [11]),
    .Q_N(_1402_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [11]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[12]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [12]),
    .Q_N(_1403_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [12]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[13]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [13]),
    .Q_N(_1404_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [13]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[14]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [14]),
    .Q_N(_1405_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [14]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[15]_reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [15]),
    .Q_N(_1406_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [15]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[16]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [16]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [16]),
    .Q_N(_1407_),
    .CLK(clknet_leaf_17_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[17]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [17]),
    .Q_N(_1408_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[18]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [18]),
    .Q_N(_1409_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[19]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [19]),
    .Q_N(_1410_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[1]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [1]),
    .Q_N(_1411_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[20]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [20]),
    .Q_N(_1412_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[21]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [21]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [21]),
    .Q_N(_1413_),
    .CLK(clknet_leaf_11_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[22]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [22]),
    .Q_N(_1414_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[23]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [23]),
    .Q_N(_1415_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[24]_reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [24]),
    .Q_N(_1416_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[25]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [25]),
    .Q_N(_1417_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[26]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [26]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [26]),
    .Q_N(_1418_),
    .CLK(clknet_leaf_10_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[27]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [27]),
    .Q_N(_1419_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[28]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [28]),
    .Q_N(_1420_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[29]_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [29]),
    .Q_N(_1421_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[2]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [2]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [2]),
    .Q_N(_1422_),
    .CLK(clknet_leaf_11_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[30]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [30]),
    .Q_N(_1423_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[31]_reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [31]),
    .Q_N(_1424_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[3]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [3]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [3]),
    .Q_N(_1425_),
    .CLK(clknet_leaf_11_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[4]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [4]),
    .Q_N(_1426_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[5]_reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [5]),
    .Q_N(_1427_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[6]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [6]),
    .Q_N(_1428_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \prescaler_lo_i.counter_value_o[7]_reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.s_count [7]),
    .Q_N(_1429_),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [7]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[8]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [8]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [8]),
    .Q_N(_1430_),
    .CLK(clknet_leaf_17_clk_i));
 sg13g2_dfrbp_2 \prescaler_lo_i.counter_value_o[9]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(\prescaler_lo_i.s_count [9]),
    .Q(\prescaler_lo_i.enable_count_i_$_MUX__S_31_B [9]),
    .Q_N(_1431_),
    .CLK(clknet_leaf_17_clk_i));
 sg13g2_dfrbp_1 \prescaler_lo_i.target_reached_o_reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(\prescaler_lo_i.target_reached_o_reg_D ),
    .Q_N(_1432_),
    .Q(\prescaler_lo_i.target_reached_o ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \r_id_o[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(id_i[0]),
    .Q(r_id_o[0]),
    .Q_N(_1433_),
    .CLK(clknet_leaf_38_clk_i));
 sg13g2_dfrbp_2 \r_id_o[1]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(id_i[1]),
    .Q(r_id_o[1]),
    .Q_N(_1434_),
    .CLK(clknet_leaf_29_clk_i));
 sg13g2_dfrbp_2 \r_id_o[2]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(id_i[2]),
    .Q(r_id_o[2]),
    .Q_N(_1435_),
    .CLK(clknet_leaf_37_clk_i));
 sg13g2_dfrbp_2 \r_id_o[3]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(id_i[3]),
    .Q(r_id_o[3]),
    .Q_N(_1436_),
    .CLK(clknet_leaf_38_clk_i));
 sg13g2_dfrbp_2 \r_id_o[4]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(id_i[4]),
    .Q(r_id_o[4]),
    .Q_N(_1437_),
    .CLK(clknet_leaf_38_clk_i));
 sg13g2_dfrbp_2 r_valid_o_reg (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(req_i),
    .Q(r_valid_o),
    .Q_N(_1438_),
    .CLK(clknet_leaf_23_clk_i));
 sg13g2_dfrbp_1 \s_addr[0]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(addr_i[0]),
    .Q_N(_1439_),
    .Q(s_addr[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_addr[1]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(addr_i[1]),
    .Q_N(_1440_),
    .Q(s_addr[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_addr[2]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(addr_i[2]),
    .Q_N(\s_addr_$_NOT__A_2_Y ),
    .Q(s_addr[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_addr[3]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(addr_i[3]),
    .Q_N(\s_addr_$_NOT__A_Y ),
    .Q(s_addr[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \s_addr[4]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(addr_i[4]),
    .Q(s_addr[4]),
    .Q_N(\s_addr_$_NOT__A_1_Y ),
    .CLK(clknet_leaf_16_clk_i));
 sg13g2_dfrbp_1 \s_addr[5]_reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(rst_ni),
    .D(addr_i[5]),
    .Q_N(_1441_),
    .Q(s_addr[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[0]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(s_cfg_hi[0]),
    .Q_N(_1255_),
    .Q(s_cfg_hi_reg[0]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[16]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0080_),
    .Q_N(_1254_),
    .Q(s_cfg_hi_reg[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[17]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0081_),
    .Q_N(_1253_),
    .Q(s_cfg_hi_reg[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[18]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0082_),
    .Q_N(_1252_),
    .Q(s_cfg_hi_reg[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[19]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0083_),
    .Q_N(_1251_),
    .Q(s_cfg_hi_reg[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[1]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0084_),
    .Q_N(_1250_),
    .Q(s_cfg_hi_reg[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[20]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0085_),
    .Q_N(_1249_),
    .Q(s_cfg_hi_reg[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[21]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0086_),
    .Q_N(_1248_),
    .Q(s_cfg_hi_reg[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[22]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0087_),
    .Q_N(_1247_),
    .Q(s_cfg_hi_reg[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[23]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0088_),
    .Q_N(_1246_),
    .Q(s_cfg_hi_reg[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[24]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0089_),
    .Q_N(_1245_),
    .Q(s_cfg_hi_reg[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[25]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0090_),
    .Q_N(_1244_),
    .Q(s_cfg_hi_reg[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[26]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0091_),
    .Q_N(_1243_),
    .Q(s_cfg_hi_reg[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[27]_reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(rst_ni),
    .D(_0092_),
    .Q_N(_1242_),
    .Q(s_cfg_hi_reg[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[28]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0093_),
    .Q_N(_1241_),
    .Q(s_cfg_hi_reg[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[29]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0094_),
    .Q_N(_1240_),
    .Q(s_cfg_hi_reg[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[2]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0095_),
    .Q_N(_1239_),
    .Q(s_cfg_hi_reg[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[30]_reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(rst_ni),
    .D(_0096_),
    .Q_N(_1238_),
    .Q(s_cfg_hi_reg[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[31]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0097_),
    .Q_N(\s_cfg_hi_$_OR__Y_A_$_MUX__Y_S_$_AND__Y_A_$_AND__Y_A ),
    .Q(s_cfg_hi_reg[31]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[3]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(s_cfg_hi[3]),
    .Q_N(_1237_),
    .Q(s_cfg_hi_reg[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[4]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0098_),
    .Q_N(_1442_),
    .Q(s_cfg_hi_reg[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[5]_reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(rst_ni),
    .D(s_cfg_hi[5]),
    .Q_N(_1236_),
    .Q(s_cfg_hi_reg[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_hi_reg[6]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0099_),
    .Q_N(\prescaler_hi_i.target_reached_o_$_MUX__A_S_$_AND__Y_A ),
    .Q(s_cfg_hi_reg[6]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \s_cfg_hi_reg[7]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0100_),
    .Q(s_cfg_hi_reg[7]),
    .Q_N(\prescaler_hi_i.enable_count_i_$_AND__Y_B_$_MUX__Y_S_$_AND__Y_B ),
    .CLK(clknet_leaf_8_clk_i));
 sg13g2_dfrbp_2 \s_cfg_lo_reg[0]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(s_cfg_lo[0]),
    .Q(s_cfg_lo_reg[0]),
    .Q_N(_1235_),
    .CLK(clknet_leaf_7_clk_i));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[16]_reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(rst_ni),
    .D(_0101_),
    .Q_N(_1234_),
    .Q(s_cfg_lo_reg[16]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[17]_reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(rst_ni),
    .D(_0102_),
    .Q_N(_1233_),
    .Q(s_cfg_lo_reg[17]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[18]_reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(rst_ni),
    .D(_0103_),
    .Q_N(_1232_),
    .Q(s_cfg_lo_reg[18]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[19]_reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(rst_ni),
    .D(_0104_),
    .Q_N(_1231_),
    .Q(s_cfg_lo_reg[19]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[1]_reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(_0105_),
    .Q_N(_1230_),
    .Q(s_cfg_lo_reg[1]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[20]_reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(rst_ni),
    .D(_0106_),
    .Q_N(_1229_),
    .Q(s_cfg_lo_reg[20]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[21]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0107_),
    .Q_N(_1228_),
    .Q(s_cfg_lo_reg[21]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[22]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0108_),
    .Q_N(_1227_),
    .Q(s_cfg_lo_reg[22]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[23]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0109_),
    .Q_N(_1226_),
    .Q(s_cfg_lo_reg[23]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[24]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0110_),
    .Q_N(_1225_),
    .Q(s_cfg_lo_reg[24]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[25]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0111_),
    .Q_N(_1224_),
    .Q(s_cfg_lo_reg[25]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[26]_reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(rst_ni),
    .D(_0112_),
    .Q_N(_1223_),
    .Q(s_cfg_lo_reg[26]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[27]_reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(rst_ni),
    .D(_0113_),
    .Q_N(_1222_),
    .Q(s_cfg_lo_reg[27]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[28]_reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(rst_ni),
    .D(_0114_),
    .Q_N(_1221_),
    .Q(s_cfg_lo_reg[28]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[29]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0115_),
    .Q_N(_1220_),
    .Q(s_cfg_lo_reg[29]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[2]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(_0116_),
    .Q_N(_1219_),
    .Q(s_cfg_lo_reg[2]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[30]_reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(rst_ni),
    .D(_0117_),
    .Q_N(_1218_),
    .Q(s_cfg_lo_reg[30]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \s_cfg_lo_reg[31]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0118_),
    .Q(s_cfg_lo_reg[31]),
    .Q_N(_1443_),
    .CLK(clknet_leaf_2_clk_i));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[3]_reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(rst_ni),
    .D(s_cfg_lo[3]),
    .Q_N(_1217_),
    .Q(s_cfg_lo_reg[3]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[4]_reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(rst_ni),
    .D(_0119_),
    .Q_N(_1444_),
    .Q(s_cfg_lo_reg[4]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 \s_cfg_lo_reg[5]_reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(rst_ni),
    .D(s_cfg_lo[5]),
    .Q_N(_1216_),
    .Q(s_cfg_lo_reg[5]),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_2 \s_cfg_lo_reg[6]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0120_),
    .Q(s_cfg_lo_reg[6]),
    .Q_N(\s_ref_clk_edge_del_$_MUX__B_S_$_AND__Y_A ),
    .CLK(clknet_leaf_8_clk_i));
 sg13g2_dfrbp_2 \s_cfg_lo_reg[7]_reg  (.RESET_B(rst_ni),
    .VSS(VSS),
    .VDD(VDD),
    .D(_0121_),
    .Q(s_cfg_lo_reg[7]),
    .Q_N(\counter_lo_i.enable_count_i_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_B ),
    .CLK(clknet_leaf_8_clk_i));
 sg13g2_dfrbp_1 s_ref_clk0_reg (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(ref_clk_i),
    .Q_N(_1445_),
    .Q(s_ref_clk0),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 s_ref_clk1_reg (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(rst_ni),
    .D(net113),
    .Q_N(_1446_),
    .Q(s_ref_clk1),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 s_ref_clk2_reg (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(net115),
    .Q_N(\s_ref_clk_edge_$_AND__Y_B ),
    .Q(s_ref_clk2),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 s_ref_clk3_reg (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(rst_ni),
    .D(net114),
    .Q_N(\s_ref_clk_edge_del_$_AND__Y_B ),
    .Q(s_ref_clk3),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbp_1 s_wen_reg (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(rst_ni),
    .D(wen_i),
    .Q_N(_1215_),
    .Q(s_wen),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo timer_unit_1 (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net1));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net92),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_0467_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout93 (.A(net97),
    .X(net93),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout94 (.A(net97),
    .X(net94),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout95 (.A(net97),
    .X(net95),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(net96),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout97 (.A(_0275_),
    .X(net97),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(net100),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net100),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout100 (.A(_0230_),
    .X(net100),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(_0230_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_0230_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_1032_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout105 (.A(_1020_),
    .X(net105),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_1009_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net111),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net111),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(net110),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net111),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_0942_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 fanout112 (.A(\counter_hi_i.enable_count_i_$_MUX__S_31_B [9]),
    .X(net112),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_0_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_1_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_1_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_2_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_2_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_3_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_3_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_4_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_4_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_5_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_5_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_6_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_6_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_7_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_7_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_8_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_8_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_9_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_9_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_10_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_10_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_11_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_11_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_12_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_12_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_13_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_13_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_14_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_14_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_15_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_15_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_16_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_16_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_17_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_17_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_18_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_18_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_19_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_19_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_20_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_20_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_21_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_21_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_22_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_22_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_23_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_23_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_24_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_24_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_25_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_25_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_26_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_26_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_27_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_27_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_28_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_28_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_29_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_29_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_30_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_30_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_31_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_31_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_32_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_32_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_33_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_33_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_34_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_34_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_35_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_35_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_36_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_36_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_37_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_37_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_leaf_38_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_38_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_0__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_1__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_2__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_3__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_4__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_4__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_5__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_5__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_6__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_6__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkbuf_3_7__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload0 (.A(clknet_3_7__leaf_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload1 (.A(clknet_leaf_0_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload2 (.A(clknet_leaf_1_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload3 (.A(clknet_leaf_2_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_37_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload5 (.A(clknet_leaf_4_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_34_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload7 (.VDD(VDD),
    .A(clknet_leaf_35_clk_i),
    .VSS(VSS));
 sg13g2_inv_1 clkload8 (.VDD(VDD),
    .A(clknet_leaf_36_clk_i),
    .VSS(VSS));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_6_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload10 (.A(clknet_leaf_7_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 clkload11 (.A(clknet_leaf_9_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_10_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_5_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload14 (.A(clknet_leaf_12_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload15 (.A(clknet_leaf_13_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_4 clkload16 (.A(clknet_leaf_14_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_25_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload18 (.VDD(VDD),
    .A(clknet_leaf_31_clk_i),
    .VSS(VSS));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_32_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_33_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload21 (.A(clknet_leaf_26_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload22 (.A(clknet_leaf_27_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload23 (.A(clknet_leaf_28_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_30_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload25 (.A(clknet_leaf_15_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload26 (.A(clknet_leaf_16_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload27 (.A(clknet_leaf_18_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_2 clkload28 (.A(clknet_leaf_23_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_inv_1 clkload29 (.VDD(VDD),
    .A(clknet_leaf_19_clk_i),
    .VSS(VSS));
 sg13g2_buf_2 clkload30 (.A(clknet_leaf_20_clk_i),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd3_1 hold113 (.A(s_ref_clk0),
    .VDD(VDD),
    .VSS(VSS),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold114 (.A(s_ref_clk2),
    .VDD(VDD),
    .VSS(VSS),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold115 (.A(s_ref_clk1),
    .VDD(VDD),
    .VSS(VSS),
    .X(net115));
 sg13g2_antennanp ANTENNA_1 (.VDD(VDD),
    .VSS(VSS),
    .A(event_lo_i));
 sg13g2_antennanp ANTENNA_2 (.VDD(VDD),
    .VSS(VSS),
    .A(id_i[0]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VDD),
    .VSS(VSS),
    .A(id_i[3]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VDD),
    .VSS(VSS),
    .A(ref_clk_i));
 sg13g2_antennanp ANTENNA_5 (.VDD(VDD),
    .VSS(VSS),
    .A(ref_clk_i));
 sg13g2_antennanp ANTENNA_6 (.VDD(VDD),
    .VSS(VSS),
    .A(id_i[0]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VDD),
    .VSS(VSS),
    .A(id_i[3]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VDD),
    .VSS(VSS),
    .A(ref_clk_i));
 sg13g2_antennanp ANTENNA_9 (.VDD(VDD),
    .VSS(VSS),
    .A(ref_clk_i));
 sg13g2_antennanp ANTENNA_10 (.VDD(VDD),
    .VSS(VSS),
    .A(id_i[0]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VDD),
    .VSS(VSS),
    .A(id_i[3]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VDD),
    .VSS(VSS),
    .A(ref_clk_i));
 sg13g2_antennanp ANTENNA_13 (.VDD(VDD),
    .VSS(VSS),
    .A(ref_clk_i));
 assign gnt_o = net2;
 assign r_opc_o = net1;
endmodule
